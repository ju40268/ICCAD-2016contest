module multiplier ( A, B, Y );
  input [15:0] A;
  input [15:0] B;
  output [31:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624;

  OR2X4 U3 ( .A(n3), .B(n4), .Y(Y[9]) );
  AND2X4 U4 ( .A(n5), .B(n6), .Y(n4) );
  AND2X4 U5 ( .A(n7), .B(n8), .Y(n6) );
  OR2X4 U6 ( .A(n9), .B(n10), .Y(n8) );
  INVX4 U7 ( .A(n11), .Y(n5) );
  AND2X4 U8 ( .A(n12), .B(n11), .Y(n3) );
  OR2X4 U9 ( .A(n13), .B(n14), .Y(n12) );
  AND2X4 U10 ( .A(n9), .B(n10), .Y(n13) );
  INVX4 U11 ( .A(n15), .Y(n10) );
  INVX4 U12 ( .A(n16), .Y(n9) );
  OR2X4 U13 ( .A(n17), .B(n18), .Y(Y[8]) );
  AND2X4 U14 ( .A(n19), .B(n20), .Y(n18) );
  AND2X4 U15 ( .A(n21), .B(n22), .Y(n20) );
  OR2X4 U16 ( .A(n23), .B(n24), .Y(n21) );
  INVX4 U17 ( .A(n25), .Y(n19) );
  AND2X4 U18 ( .A(n26), .B(n25), .Y(n17) );
  OR2X4 U19 ( .A(n27), .B(n28), .Y(n26) );
  AND2X4 U20 ( .A(n23), .B(n24), .Y(n27) );
  INVX4 U21 ( .A(n29), .Y(n24) );
  INVX4 U22 ( .A(n30), .Y(n23) );
  OR2X4 U23 ( .A(n31), .B(n32), .Y(Y[7]) );
  AND2X4 U24 ( .A(n33), .B(n34), .Y(n32) );
  AND2X4 U25 ( .A(n35), .B(n36), .Y(n34) );
  OR2X4 U26 ( .A(n37), .B(n38), .Y(n35) );
  INVX4 U27 ( .A(n39), .Y(n33) );
  AND2X4 U28 ( .A(n40), .B(n39), .Y(n31) );
  OR2X4 U29 ( .A(n41), .B(n42), .Y(n40) );
  AND2X4 U30 ( .A(n37), .B(n38), .Y(n41) );
  INVX4 U31 ( .A(n43), .Y(n38) );
  INVX4 U32 ( .A(n44), .Y(n37) );
  OR2X4 U33 ( .A(n45), .B(n46), .Y(Y[6]) );
  AND2X4 U34 ( .A(n47), .B(n48), .Y(n46) );
  AND2X4 U35 ( .A(n49), .B(n50), .Y(n48) );
  OR2X4 U36 ( .A(n51), .B(n52), .Y(n49) );
  INVX4 U37 ( .A(n53), .Y(n47) );
  AND2X4 U38 ( .A(n54), .B(n53), .Y(n45) );
  OR2X4 U39 ( .A(n55), .B(n56), .Y(n54) );
  AND2X4 U40 ( .A(n51), .B(n52), .Y(n55) );
  INVX4 U41 ( .A(n57), .Y(n52) );
  INVX4 U42 ( .A(n58), .Y(n51) );
  OR2X4 U43 ( .A(n59), .B(n60), .Y(Y[5]) );
  AND2X4 U44 ( .A(n61), .B(n62), .Y(n60) );
  AND2X4 U45 ( .A(n63), .B(n64), .Y(n62) );
  OR2X4 U46 ( .A(n65), .B(n66), .Y(n63) );
  INVX4 U47 ( .A(n67), .Y(n61) );
  AND2X4 U48 ( .A(n68), .B(n67), .Y(n59) );
  OR2X4 U49 ( .A(n69), .B(n70), .Y(n68) );
  AND2X4 U50 ( .A(n65), .B(n66), .Y(n69) );
  INVX4 U51 ( .A(n71), .Y(n66) );
  INVX4 U52 ( .A(n72), .Y(n65) );
  OR2X4 U53 ( .A(n73), .B(n74), .Y(Y[4]) );
  AND2X4 U54 ( .A(n75), .B(n76), .Y(n74) );
  AND2X4 U55 ( .A(n77), .B(n78), .Y(n76) );
  OR2X4 U56 ( .A(n79), .B(n80), .Y(n77) );
  INVX4 U57 ( .A(n81), .Y(n75) );
  AND2X4 U58 ( .A(n82), .B(n81), .Y(n73) );
  OR2X4 U59 ( .A(n83), .B(n84), .Y(n82) );
  AND2X4 U60 ( .A(n79), .B(n80), .Y(n83) );
  INVX4 U61 ( .A(n85), .Y(n80) );
  INVX4 U62 ( .A(n86), .Y(n79) );
  OR2X4 U63 ( .A(n87), .B(n88), .Y(Y[3]) );
  AND2X4 U64 ( .A(n89), .B(n90), .Y(n88) );
  AND2X4 U65 ( .A(n91), .B(n92), .Y(n90) );
  OR2X4 U66 ( .A(n93), .B(n94), .Y(n91) );
  INVX4 U67 ( .A(n95), .Y(n89) );
  AND2X4 U68 ( .A(n95), .B(n96), .Y(n87) );
  OR2X4 U69 ( .A(n97), .B(n98), .Y(n96) );
  AND2X4 U70 ( .A(n93), .B(n94), .Y(n97) );
  INVX4 U71 ( .A(n99), .Y(n94) );
  INVX4 U72 ( .A(n100), .Y(n93) );
  OR2X4 U73 ( .A(n101), .B(n102), .Y(Y[31]) );
  OR2X4 U74 ( .A(n103), .B(n104), .Y(n102) );
  AND2X4 U75 ( .A(n105), .B(n106), .Y(n104) );
  AND2X4 U76 ( .A(n106), .B(n107), .Y(n103) );
  OR2X4 U77 ( .A(n108), .B(n109), .Y(n101) );
  AND2X4 U78 ( .A(A[15]), .B(n110), .Y(n109) );
  OR2X4 U79 ( .A(n111), .B(n112), .Y(Y[30]) );
  AND2X4 U80 ( .A(n113), .B(n106), .Y(n112) );
  NOR2X4 U81 ( .A(n106), .B(n113), .Y(n111) );
  NOR2X4 U82 ( .A(n105), .B(n107), .Y(n113) );
  NAND2X4 U83 ( .A(n114), .B(n115), .Y(n107) );
  OR2X4 U84 ( .A(n116), .B(n117), .Y(n106) );
  AND2X4 U85 ( .A(n118), .B(n110), .Y(n117) );
  AND2X4 U86 ( .A(n119), .B(n120), .Y(n116) );
  AND2X4 U87 ( .A(A[15]), .B(n121), .Y(n120) );
  AND2X4 U88 ( .A(n122), .B(B[15]), .Y(n119) );
  OR2X4 U89 ( .A(n123), .B(n124), .Y(Y[2]) );
  OR2X4 U90 ( .A(n125), .B(n126), .Y(n124) );
  AND2X4 U91 ( .A(n127), .B(n128), .Y(n126) );
  AND2X4 U92 ( .A(B[0]), .B(n129), .Y(n127) );
  OR2X4 U93 ( .A(n130), .B(n131), .Y(n129) );
  AND2X4 U94 ( .A(A[2]), .B(n132), .Y(n130) );
  AND2X4 U95 ( .A(n133), .B(n134), .Y(n125) );
  OR2X4 U96 ( .A(n135), .B(n136), .Y(n133) );
  OR2X4 U97 ( .A(n137), .B(n138), .Y(n136) );
  OR2X4 U98 ( .A(n139), .B(n140), .Y(n135) );
  AND2X4 U99 ( .A(n141), .B(B[1]), .Y(n140) );
  AND2X4 U100 ( .A(n142), .B(n132), .Y(n139) );
  AND2X4 U101 ( .A(n143), .B(n144), .Y(n123) );
  AND2X4 U102 ( .A(Y[0]), .B(n145), .Y(n143) );
  AND2X4 U103 ( .A(n146), .B(n115), .Y(Y[29]) );
  OR2X4 U104 ( .A(n147), .B(n148), .Y(n115) );
  OR2X4 U105 ( .A(n105), .B(n149), .Y(n148) );
  AND2X4 U106 ( .A(n150), .B(n151), .Y(n149) );
  NOR2X4 U107 ( .A(n150), .B(n151), .Y(n105) );
  INVX4 U108 ( .A(n152), .Y(n150) );
  AND2X4 U109 ( .A(n153), .B(n154), .Y(n147) );
  OR2X4 U110 ( .A(n155), .B(n156), .Y(n153) );
  OR2X4 U111 ( .A(n157), .B(n158), .Y(n146) );
  OR2X4 U112 ( .A(n159), .B(n160), .Y(n158) );
  AND2X4 U113 ( .A(n161), .B(n114), .Y(n160) );
  NAND2X4 U114 ( .A(n162), .B(n163), .Y(n114) );
  OR2X4 U115 ( .A(n163), .B(n162), .Y(n161) );
  OR2X4 U116 ( .A(n164), .B(n165), .Y(n162) );
  AND2X4 U117 ( .A(n151), .B(n152), .Y(n165) );
  NOR2X4 U118 ( .A(n151), .B(n152), .Y(n164) );
  OR2X4 U119 ( .A(n166), .B(n167), .Y(n152) );
  AND2X4 U120 ( .A(n168), .B(n169), .Y(n166) );
  OR2X4 U121 ( .A(n170), .B(n171), .Y(n151) );
  AND2X4 U122 ( .A(n172), .B(n110), .Y(n171) );
  OR2X4 U123 ( .A(n118), .B(n173), .Y(n172) );
  AND2X4 U124 ( .A(A[15]), .B(n174), .Y(n173) );
  AND2X4 U125 ( .A(n175), .B(A[14]), .Y(n118) );
  AND2X4 U126 ( .A(n122), .B(n176), .Y(n170) );
  OR2X4 U127 ( .A(n177), .B(n178), .Y(n176) );
  OR2X4 U128 ( .A(n179), .B(n180), .Y(n178) );
  AND2X4 U129 ( .A(n181), .B(n175), .Y(n180) );
  OR2X4 U130 ( .A(n174), .B(n182), .Y(n181) );
  AND2X4 U131 ( .A(n174), .B(n183), .Y(n179) );
  INVX4 U132 ( .A(A[14]), .Y(n174) );
  OR2X4 U133 ( .A(n184), .B(n108), .Y(n177) );
  AND2X4 U134 ( .A(n185), .B(B[15]), .Y(n108) );
  AND2X4 U135 ( .A(A[15]), .B(n186), .Y(n185) );
  AND2X4 U136 ( .A(n183), .B(n182), .Y(n184) );
  INVX4 U137 ( .A(n110), .Y(n122) );
  OR2X4 U138 ( .A(n187), .B(n188), .Y(n110) );
  AND2X4 U139 ( .A(n189), .B(n190), .Y(n187) );
  OR2X4 U140 ( .A(n191), .B(n186), .Y(n189) );
  NOR2X4 U141 ( .A(n155), .B(n156), .Y(n157) );
  AND2X4 U142 ( .A(n192), .B(n193), .Y(Y[28]) );
  NAND2X4 U143 ( .A(n194), .B(n156), .Y(n193) );
  OR2X4 U144 ( .A(n156), .B(n194), .Y(n192) );
  OR2X4 U145 ( .A(n155), .B(n159), .Y(n194) );
  INVX4 U146 ( .A(n154), .Y(n159) );
  OR2X4 U147 ( .A(n195), .B(n196), .Y(n154) );
  OR2X4 U148 ( .A(n197), .B(n198), .Y(n196) );
  AND2X4 U149 ( .A(n199), .B(n198), .Y(n155) );
  OR2X4 U150 ( .A(n200), .B(n163), .Y(n198) );
  NOR2X4 U151 ( .A(n201), .B(n202), .Y(n163) );
  AND2X4 U152 ( .A(n201), .B(n202), .Y(n200) );
  NOR2X4 U153 ( .A(n203), .B(n204), .Y(n202) );
  AND2X4 U154 ( .A(n205), .B(n206), .Y(n204) );
  AND2X4 U155 ( .A(n207), .B(n169), .Y(n206) );
  OR2X4 U156 ( .A(n208), .B(n209), .Y(n169) );
  OR2X4 U157 ( .A(n210), .B(n211), .Y(n207) );
  INVX4 U158 ( .A(n168), .Y(n205) );
  AND2X4 U159 ( .A(n168), .B(n212), .Y(n203) );
  OR2X4 U160 ( .A(n213), .B(n167), .Y(n212) );
  AND2X4 U161 ( .A(n209), .B(n208), .Y(n167) );
  AND2X4 U162 ( .A(n210), .B(n211), .Y(n213) );
  INVX4 U163 ( .A(n208), .Y(n211) );
  AND2X4 U164 ( .A(A[15]), .B(B[13]), .Y(n208) );
  INVX4 U165 ( .A(n209), .Y(n210) );
  OR2X4 U166 ( .A(n214), .B(n215), .Y(n209) );
  AND2X4 U167 ( .A(n216), .B(n217), .Y(n214) );
  OR2X4 U168 ( .A(n218), .B(n219), .Y(n168) );
  AND2X4 U169 ( .A(n220), .B(n221), .Y(n219) );
  OR2X4 U170 ( .A(n222), .B(n223), .Y(n221) );
  AND2X4 U171 ( .A(n191), .B(n121), .Y(n223) );
  AND2X4 U172 ( .A(n186), .B(n224), .Y(n222) );
  INVX4 U173 ( .A(n190), .Y(n220) );
  AND2X4 U174 ( .A(n225), .B(n190), .Y(n218) );
  OR2X4 U175 ( .A(n226), .B(n227), .Y(n190) );
  AND2X4 U176 ( .A(n228), .B(n229), .Y(n226) );
  OR2X4 U177 ( .A(A[12]), .B(A[13]), .Y(n228) );
  OR2X4 U178 ( .A(n230), .B(n188), .Y(n225) );
  AND2X4 U179 ( .A(n186), .B(n191), .Y(n188) );
  AND2X4 U180 ( .A(n224), .B(n121), .Y(n230) );
  INVX4 U181 ( .A(n186), .Y(n121) );
  AND2X4 U182 ( .A(A[14]), .B(B[14]), .Y(n186) );
  INVX4 U183 ( .A(n191), .Y(n224) );
  AND2X4 U184 ( .A(B[15]), .B(A[13]), .Y(n191) );
  NOR2X4 U185 ( .A(n231), .B(n232), .Y(n201) );
  OR2X4 U186 ( .A(n233), .B(n234), .Y(n232) );
  AND2X4 U187 ( .A(n235), .B(n236), .Y(n231) );
  OR2X4 U188 ( .A(n195), .B(n197), .Y(n199) );
  AND2X4 U189 ( .A(n237), .B(n238), .Y(n156) );
  AND2X4 U190 ( .A(n239), .B(n238), .Y(Y[27]) );
  OR2X4 U191 ( .A(n240), .B(n241), .Y(n238) );
  AND2X4 U192 ( .A(n242), .B(n243), .Y(n240) );
  OR2X4 U193 ( .A(n244), .B(n245), .Y(n242) );
  OR2X4 U194 ( .A(n246), .B(n247), .Y(n239) );
  OR2X4 U195 ( .A(n248), .B(n249), .Y(n247) );
  AND2X4 U196 ( .A(n250), .B(n237), .Y(n249) );
  NAND2X4 U197 ( .A(n251), .B(n252), .Y(n237) );
  OR2X4 U198 ( .A(n252), .B(n251), .Y(n250) );
  INVX4 U199 ( .A(n241), .Y(n251) );
  OR2X4 U200 ( .A(n253), .B(n254), .Y(n241) );
  NOR2X4 U201 ( .A(n195), .B(n197), .Y(n254) );
  AND2X4 U202 ( .A(n197), .B(n195), .Y(n253) );
  OR2X4 U203 ( .A(n255), .B(n256), .Y(n195) );
  OR2X4 U204 ( .A(n257), .B(n258), .Y(n256) );
  AND2X4 U205 ( .A(n259), .B(n260), .Y(n258) );
  OR2X4 U206 ( .A(n261), .B(n233), .Y(n260) );
  NOR2X4 U207 ( .A(n262), .B(n263), .Y(n233) );
  AND2X4 U208 ( .A(n262), .B(n263), .Y(n261) );
  AND2X4 U209 ( .A(n264), .B(n235), .Y(n257) );
  AND2X4 U210 ( .A(n263), .B(n236), .Y(n264) );
  AND2X4 U211 ( .A(n234), .B(n262), .Y(n255) );
  INVX4 U212 ( .A(n236), .Y(n262) );
  OR2X4 U213 ( .A(n265), .B(n266), .Y(n236) );
  AND2X4 U214 ( .A(n267), .B(n268), .Y(n265) );
  NOR2X4 U215 ( .A(n259), .B(n263), .Y(n234) );
  OR2X4 U216 ( .A(n175), .B(n269), .Y(n263) );
  INVX4 U217 ( .A(n235), .Y(n259) );
  OR2X4 U218 ( .A(n270), .B(n271), .Y(n235) );
  AND2X4 U219 ( .A(n272), .B(n273), .Y(n271) );
  AND2X4 U220 ( .A(n274), .B(n217), .Y(n273) );
  OR2X4 U221 ( .A(n275), .B(n276), .Y(n217) );
  OR2X4 U222 ( .A(n277), .B(n278), .Y(n274) );
  INVX4 U223 ( .A(n216), .Y(n272) );
  AND2X4 U224 ( .A(n216), .B(n279), .Y(n270) );
  OR2X4 U225 ( .A(n280), .B(n215), .Y(n279) );
  AND2X4 U226 ( .A(n276), .B(n275), .Y(n215) );
  AND2X4 U227 ( .A(n277), .B(n278), .Y(n280) );
  INVX4 U228 ( .A(n275), .Y(n278) );
  AND2X4 U229 ( .A(A[14]), .B(B[13]), .Y(n275) );
  INVX4 U230 ( .A(n276), .Y(n277) );
  OR2X4 U231 ( .A(n281), .B(n282), .Y(n276) );
  AND2X4 U232 ( .A(n283), .B(n284), .Y(n281) );
  OR2X4 U233 ( .A(n285), .B(n286), .Y(n216) );
  AND2X4 U234 ( .A(n287), .B(n288), .Y(n286) );
  OR2X4 U235 ( .A(n289), .B(n290), .Y(n288) );
  AND2X4 U236 ( .A(A[13]), .B(n291), .Y(n290) );
  OR2X4 U237 ( .A(n292), .B(n293), .Y(n291) );
  AND2X4 U238 ( .A(B[14]), .B(n294), .Y(n292) );
  AND2X4 U239 ( .A(A[12]), .B(n295), .Y(n289) );
  OR2X4 U240 ( .A(n296), .B(n297), .Y(n295) );
  AND2X4 U241 ( .A(B[15]), .B(n298), .Y(n296) );
  INVX4 U242 ( .A(n229), .Y(n287) );
  AND2X4 U243 ( .A(n299), .B(n229), .Y(n285) );
  OR2X4 U244 ( .A(n300), .B(n301), .Y(n229) );
  AND2X4 U245 ( .A(n302), .B(n303), .Y(n300) );
  OR2X4 U246 ( .A(A[11]), .B(A[12]), .Y(n302) );
  OR2X4 U247 ( .A(n227), .B(n304), .Y(n299) );
  AND2X4 U248 ( .A(n294), .B(n298), .Y(n304) );
  INVX4 U249 ( .A(A[13]), .Y(n298) );
  AND2X4 U250 ( .A(n305), .B(A[13]), .Y(n227) );
  AND2X4 U251 ( .A(A[12]), .B(n306), .Y(n305) );
  NOR2X4 U252 ( .A(n307), .B(n308), .Y(n197) );
  AND2X4 U253 ( .A(n309), .B(n310), .Y(n307) );
  NOR2X4 U254 ( .A(n244), .B(n245), .Y(n246) );
  AND2X4 U255 ( .A(n311), .B(n312), .Y(Y[26]) );
  NAND2X4 U256 ( .A(n313), .B(n245), .Y(n312) );
  OR2X4 U257 ( .A(n245), .B(n313), .Y(n311) );
  OR2X4 U258 ( .A(n244), .B(n248), .Y(n313) );
  INVX4 U259 ( .A(n243), .Y(n248) );
  OR2X4 U260 ( .A(n314), .B(n315), .Y(n243) );
  OR2X4 U261 ( .A(n316), .B(n317), .Y(n315) );
  AND2X4 U262 ( .A(n318), .B(n317), .Y(n244) );
  OR2X4 U263 ( .A(n319), .B(n252), .Y(n317) );
  NOR2X4 U264 ( .A(n320), .B(n321), .Y(n252) );
  AND2X4 U265 ( .A(n320), .B(n321), .Y(n319) );
  NOR2X4 U266 ( .A(n322), .B(n323), .Y(n321) );
  AND2X4 U267 ( .A(n324), .B(n325), .Y(n323) );
  AND2X4 U268 ( .A(n326), .B(n310), .Y(n325) );
  OR2X4 U269 ( .A(n327), .B(n328), .Y(n310) );
  OR2X4 U270 ( .A(n329), .B(n330), .Y(n326) );
  INVX4 U271 ( .A(n309), .Y(n324) );
  AND2X4 U272 ( .A(n309), .B(n331), .Y(n322) );
  OR2X4 U273 ( .A(n332), .B(n308), .Y(n331) );
  AND2X4 U274 ( .A(n328), .B(n327), .Y(n308) );
  AND2X4 U275 ( .A(n329), .B(n330), .Y(n332) );
  INVX4 U276 ( .A(n327), .Y(n330) );
  AND2X4 U277 ( .A(A[15]), .B(B[11]), .Y(n327) );
  INVX4 U278 ( .A(n328), .Y(n329) );
  OR2X4 U279 ( .A(n333), .B(n334), .Y(n328) );
  AND2X4 U280 ( .A(n335), .B(n336), .Y(n333) );
  OR2X4 U281 ( .A(n337), .B(n338), .Y(n309) );
  AND2X4 U282 ( .A(n339), .B(n340), .Y(n338) );
  AND2X4 U283 ( .A(n341), .B(n268), .Y(n340) );
  OR2X4 U284 ( .A(n342), .B(n343), .Y(n268) );
  OR2X4 U285 ( .A(n344), .B(n345), .Y(n341) );
  INVX4 U286 ( .A(n267), .Y(n339) );
  AND2X4 U287 ( .A(n267), .B(n346), .Y(n337) );
  OR2X4 U288 ( .A(n347), .B(n266), .Y(n346) );
  AND2X4 U289 ( .A(n343), .B(n342), .Y(n266) );
  AND2X4 U290 ( .A(n344), .B(n345), .Y(n347) );
  INVX4 U291 ( .A(n342), .Y(n345) );
  AND2X4 U292 ( .A(A[14]), .B(B[12]), .Y(n342) );
  INVX4 U293 ( .A(n343), .Y(n344) );
  OR2X4 U294 ( .A(n348), .B(n349), .Y(n343) );
  AND2X4 U295 ( .A(n350), .B(n351), .Y(n348) );
  OR2X4 U296 ( .A(n352), .B(n353), .Y(n267) );
  AND2X4 U297 ( .A(n354), .B(n355), .Y(n353) );
  AND2X4 U298 ( .A(n356), .B(n284), .Y(n355) );
  OR2X4 U299 ( .A(n357), .B(n358), .Y(n284) );
  OR2X4 U300 ( .A(n359), .B(n360), .Y(n356) );
  INVX4 U301 ( .A(n283), .Y(n354) );
  AND2X4 U302 ( .A(n283), .B(n361), .Y(n352) );
  OR2X4 U303 ( .A(n362), .B(n282), .Y(n361) );
  AND2X4 U304 ( .A(n358), .B(n357), .Y(n282) );
  AND2X4 U305 ( .A(n359), .B(n360), .Y(n362) );
  INVX4 U306 ( .A(n357), .Y(n360) );
  AND2X4 U307 ( .A(A[13]), .B(B[13]), .Y(n357) );
  INVX4 U308 ( .A(n358), .Y(n359) );
  OR2X4 U309 ( .A(n363), .B(n364), .Y(n358) );
  AND2X4 U310 ( .A(n365), .B(n366), .Y(n363) );
  OR2X4 U311 ( .A(n367), .B(n368), .Y(n283) );
  AND2X4 U312 ( .A(n369), .B(n370), .Y(n368) );
  OR2X4 U313 ( .A(n371), .B(n372), .Y(n370) );
  AND2X4 U314 ( .A(A[12]), .B(n373), .Y(n372) );
  OR2X4 U315 ( .A(n374), .B(n293), .Y(n373) );
  AND2X4 U316 ( .A(B[14]), .B(n375), .Y(n374) );
  AND2X4 U317 ( .A(A[11]), .B(n376), .Y(n371) );
  OR2X4 U318 ( .A(n377), .B(n297), .Y(n376) );
  AND2X4 U319 ( .A(B[15]), .B(n294), .Y(n377) );
  INVX4 U320 ( .A(n303), .Y(n369) );
  AND2X4 U321 ( .A(n378), .B(n303), .Y(n367) );
  OR2X4 U322 ( .A(n379), .B(n380), .Y(n303) );
  AND2X4 U323 ( .A(n381), .B(n382), .Y(n379) );
  OR2X4 U324 ( .A(A[10]), .B(A[11]), .Y(n381) );
  OR2X4 U325 ( .A(n301), .B(n383), .Y(n378) );
  AND2X4 U326 ( .A(n375), .B(n294), .Y(n383) );
  INVX4 U327 ( .A(A[12]), .Y(n294) );
  AND2X4 U328 ( .A(n384), .B(A[12]), .Y(n301) );
  AND2X4 U329 ( .A(A[11]), .B(n306), .Y(n384) );
  NOR2X4 U330 ( .A(n385), .B(n386), .Y(n320) );
  OR2X4 U331 ( .A(n387), .B(n388), .Y(n386) );
  AND2X4 U332 ( .A(n389), .B(n390), .Y(n385) );
  OR2X4 U333 ( .A(n314), .B(n316), .Y(n318) );
  AND2X4 U334 ( .A(n391), .B(n392), .Y(n245) );
  AND2X4 U335 ( .A(n393), .B(n392), .Y(Y[25]) );
  OR2X4 U336 ( .A(n394), .B(n395), .Y(n392) );
  AND2X4 U337 ( .A(n396), .B(n397), .Y(n394) );
  OR2X4 U338 ( .A(n398), .B(n399), .Y(n396) );
  OR2X4 U339 ( .A(n400), .B(n401), .Y(n393) );
  OR2X4 U340 ( .A(n402), .B(n403), .Y(n401) );
  AND2X4 U341 ( .A(n404), .B(n391), .Y(n403) );
  NAND2X4 U342 ( .A(n405), .B(n406), .Y(n391) );
  OR2X4 U343 ( .A(n406), .B(n405), .Y(n404) );
  INVX4 U344 ( .A(n395), .Y(n405) );
  OR2X4 U345 ( .A(n407), .B(n408), .Y(n395) );
  NOR2X4 U346 ( .A(n314), .B(n316), .Y(n408) );
  AND2X4 U347 ( .A(n316), .B(n314), .Y(n407) );
  OR2X4 U348 ( .A(n409), .B(n410), .Y(n314) );
  OR2X4 U349 ( .A(n411), .B(n412), .Y(n410) );
  AND2X4 U350 ( .A(n413), .B(n414), .Y(n412) );
  OR2X4 U351 ( .A(n415), .B(n387), .Y(n414) );
  NOR2X4 U352 ( .A(n416), .B(n417), .Y(n387) );
  AND2X4 U353 ( .A(n416), .B(n417), .Y(n415) );
  AND2X4 U354 ( .A(n418), .B(n389), .Y(n411) );
  AND2X4 U355 ( .A(n417), .B(n390), .Y(n418) );
  AND2X4 U356 ( .A(n388), .B(n416), .Y(n409) );
  INVX4 U357 ( .A(n390), .Y(n416) );
  OR2X4 U358 ( .A(n419), .B(n420), .Y(n390) );
  AND2X4 U359 ( .A(n421), .B(n422), .Y(n419) );
  NOR2X4 U360 ( .A(n413), .B(n417), .Y(n388) );
  OR2X4 U361 ( .A(n175), .B(n423), .Y(n417) );
  INVX4 U362 ( .A(n389), .Y(n413) );
  OR2X4 U363 ( .A(n424), .B(n425), .Y(n389) );
  AND2X4 U364 ( .A(n426), .B(n427), .Y(n425) );
  AND2X4 U365 ( .A(n428), .B(n336), .Y(n427) );
  OR2X4 U366 ( .A(n429), .B(n430), .Y(n336) );
  OR2X4 U367 ( .A(n431), .B(n432), .Y(n428) );
  INVX4 U368 ( .A(n335), .Y(n426) );
  AND2X4 U369 ( .A(n335), .B(n433), .Y(n424) );
  OR2X4 U370 ( .A(n434), .B(n334), .Y(n433) );
  AND2X4 U371 ( .A(n430), .B(n429), .Y(n334) );
  AND2X4 U372 ( .A(n431), .B(n432), .Y(n434) );
  INVX4 U373 ( .A(n429), .Y(n432) );
  AND2X4 U374 ( .A(A[14]), .B(B[11]), .Y(n429) );
  INVX4 U375 ( .A(n430), .Y(n431) );
  OR2X4 U376 ( .A(n435), .B(n436), .Y(n430) );
  AND2X4 U377 ( .A(n437), .B(n438), .Y(n435) );
  OR2X4 U378 ( .A(n439), .B(n440), .Y(n335) );
  AND2X4 U379 ( .A(n441), .B(n442), .Y(n440) );
  AND2X4 U380 ( .A(n443), .B(n351), .Y(n442) );
  OR2X4 U381 ( .A(n444), .B(n445), .Y(n351) );
  OR2X4 U382 ( .A(n446), .B(n447), .Y(n443) );
  INVX4 U383 ( .A(n350), .Y(n441) );
  AND2X4 U384 ( .A(n350), .B(n448), .Y(n439) );
  OR2X4 U385 ( .A(n449), .B(n349), .Y(n448) );
  AND2X4 U386 ( .A(n445), .B(n444), .Y(n349) );
  AND2X4 U387 ( .A(n446), .B(n447), .Y(n449) );
  INVX4 U388 ( .A(n444), .Y(n447) );
  AND2X4 U389 ( .A(A[13]), .B(B[12]), .Y(n444) );
  INVX4 U390 ( .A(n445), .Y(n446) );
  OR2X4 U391 ( .A(n450), .B(n451), .Y(n445) );
  AND2X4 U392 ( .A(n452), .B(n453), .Y(n450) );
  OR2X4 U393 ( .A(n454), .B(n455), .Y(n350) );
  AND2X4 U394 ( .A(n456), .B(n457), .Y(n455) );
  AND2X4 U395 ( .A(n458), .B(n366), .Y(n457) );
  OR2X4 U396 ( .A(n459), .B(n460), .Y(n366) );
  OR2X4 U397 ( .A(n461), .B(n462), .Y(n458) );
  INVX4 U398 ( .A(n365), .Y(n456) );
  AND2X4 U399 ( .A(n365), .B(n463), .Y(n454) );
  OR2X4 U400 ( .A(n464), .B(n364), .Y(n463) );
  AND2X4 U401 ( .A(n460), .B(n459), .Y(n364) );
  AND2X4 U402 ( .A(n461), .B(n462), .Y(n464) );
  INVX4 U403 ( .A(n459), .Y(n462) );
  AND2X4 U404 ( .A(A[12]), .B(B[13]), .Y(n459) );
  INVX4 U405 ( .A(n460), .Y(n461) );
  OR2X4 U406 ( .A(n465), .B(n466), .Y(n460) );
  AND2X4 U407 ( .A(n467), .B(n468), .Y(n465) );
  OR2X4 U408 ( .A(n469), .B(n470), .Y(n365) );
  AND2X4 U409 ( .A(n471), .B(n472), .Y(n470) );
  OR2X4 U410 ( .A(n473), .B(n474), .Y(n472) );
  AND2X4 U411 ( .A(A[11]), .B(n475), .Y(n474) );
  OR2X4 U412 ( .A(n476), .B(n293), .Y(n475) );
  AND2X4 U413 ( .A(B[14]), .B(n477), .Y(n476) );
  AND2X4 U414 ( .A(A[10]), .B(n478), .Y(n473) );
  OR2X4 U415 ( .A(n479), .B(n297), .Y(n478) );
  AND2X4 U416 ( .A(B[15]), .B(n375), .Y(n479) );
  INVX4 U417 ( .A(n382), .Y(n471) );
  AND2X4 U418 ( .A(n480), .B(n382), .Y(n469) );
  OR2X4 U419 ( .A(n481), .B(n482), .Y(n382) );
  AND2X4 U420 ( .A(n483), .B(n484), .Y(n481) );
  OR2X4 U421 ( .A(A[10]), .B(A[9]), .Y(n483) );
  OR2X4 U422 ( .A(n380), .B(n485), .Y(n480) );
  AND2X4 U423 ( .A(n477), .B(n375), .Y(n485) );
  INVX4 U424 ( .A(A[11]), .Y(n375) );
  AND2X4 U425 ( .A(n486), .B(A[11]), .Y(n380) );
  AND2X4 U426 ( .A(A[10]), .B(n306), .Y(n486) );
  NOR2X4 U427 ( .A(n487), .B(n488), .Y(n316) );
  AND2X4 U428 ( .A(n489), .B(n490), .Y(n487) );
  NOR2X4 U429 ( .A(n398), .B(n399), .Y(n400) );
  AND2X4 U430 ( .A(n491), .B(n492), .Y(Y[24]) );
  NAND2X4 U431 ( .A(n493), .B(n399), .Y(n492) );
  OR2X4 U432 ( .A(n399), .B(n493), .Y(n491) );
  OR2X4 U433 ( .A(n398), .B(n402), .Y(n493) );
  INVX4 U434 ( .A(n397), .Y(n402) );
  OR2X4 U435 ( .A(n494), .B(n495), .Y(n397) );
  OR2X4 U436 ( .A(n496), .B(n497), .Y(n495) );
  AND2X4 U437 ( .A(n498), .B(n497), .Y(n398) );
  OR2X4 U438 ( .A(n499), .B(n406), .Y(n497) );
  NOR2X4 U439 ( .A(n500), .B(n501), .Y(n406) );
  AND2X4 U440 ( .A(n500), .B(n501), .Y(n499) );
  NOR2X4 U441 ( .A(n502), .B(n503), .Y(n501) );
  AND2X4 U442 ( .A(n504), .B(n505), .Y(n503) );
  AND2X4 U443 ( .A(n506), .B(n490), .Y(n505) );
  OR2X4 U444 ( .A(n507), .B(n508), .Y(n490) );
  OR2X4 U445 ( .A(n509), .B(n510), .Y(n506) );
  INVX4 U446 ( .A(n489), .Y(n504) );
  AND2X4 U447 ( .A(n489), .B(n511), .Y(n502) );
  OR2X4 U448 ( .A(n512), .B(n488), .Y(n511) );
  AND2X4 U449 ( .A(n508), .B(n507), .Y(n488) );
  AND2X4 U450 ( .A(n509), .B(n510), .Y(n512) );
  INVX4 U451 ( .A(n507), .Y(n510) );
  AND2X4 U452 ( .A(B[9]), .B(A[15]), .Y(n507) );
  INVX4 U453 ( .A(n508), .Y(n509) );
  OR2X4 U454 ( .A(n513), .B(n514), .Y(n508) );
  AND2X4 U455 ( .A(n515), .B(n516), .Y(n513) );
  OR2X4 U456 ( .A(n517), .B(n518), .Y(n489) );
  AND2X4 U457 ( .A(n519), .B(n520), .Y(n518) );
  AND2X4 U458 ( .A(n521), .B(n422), .Y(n520) );
  OR2X4 U459 ( .A(n522), .B(n523), .Y(n422) );
  OR2X4 U460 ( .A(n524), .B(n525), .Y(n521) );
  INVX4 U461 ( .A(n421), .Y(n519) );
  AND2X4 U462 ( .A(n421), .B(n526), .Y(n517) );
  OR2X4 U463 ( .A(n527), .B(n420), .Y(n526) );
  AND2X4 U464 ( .A(n523), .B(n522), .Y(n420) );
  AND2X4 U465 ( .A(n524), .B(n525), .Y(n527) );
  INVX4 U466 ( .A(n522), .Y(n525) );
  AND2X4 U467 ( .A(A[14]), .B(B[10]), .Y(n522) );
  INVX4 U468 ( .A(n523), .Y(n524) );
  OR2X4 U469 ( .A(n528), .B(n529), .Y(n523) );
  AND2X4 U470 ( .A(n530), .B(n531), .Y(n528) );
  OR2X4 U471 ( .A(n532), .B(n533), .Y(n421) );
  AND2X4 U472 ( .A(n534), .B(n535), .Y(n533) );
  AND2X4 U473 ( .A(n536), .B(n438), .Y(n535) );
  OR2X4 U474 ( .A(n537), .B(n538), .Y(n438) );
  OR2X4 U475 ( .A(n539), .B(n540), .Y(n536) );
  INVX4 U476 ( .A(n437), .Y(n534) );
  AND2X4 U477 ( .A(n437), .B(n541), .Y(n532) );
  OR2X4 U478 ( .A(n542), .B(n436), .Y(n541) );
  AND2X4 U479 ( .A(n538), .B(n537), .Y(n436) );
  AND2X4 U480 ( .A(n539), .B(n540), .Y(n542) );
  INVX4 U481 ( .A(n537), .Y(n540) );
  AND2X4 U482 ( .A(A[13]), .B(B[11]), .Y(n537) );
  INVX4 U483 ( .A(n538), .Y(n539) );
  OR2X4 U484 ( .A(n543), .B(n544), .Y(n538) );
  AND2X4 U485 ( .A(n545), .B(n546), .Y(n543) );
  OR2X4 U486 ( .A(n547), .B(n548), .Y(n437) );
  AND2X4 U487 ( .A(n549), .B(n550), .Y(n548) );
  AND2X4 U488 ( .A(n551), .B(n453), .Y(n550) );
  OR2X4 U489 ( .A(n552), .B(n553), .Y(n453) );
  OR2X4 U490 ( .A(n554), .B(n555), .Y(n551) );
  INVX4 U491 ( .A(n452), .Y(n549) );
  AND2X4 U492 ( .A(n452), .B(n556), .Y(n547) );
  OR2X4 U493 ( .A(n557), .B(n451), .Y(n556) );
  AND2X4 U494 ( .A(n553), .B(n552), .Y(n451) );
  AND2X4 U495 ( .A(n554), .B(n555), .Y(n557) );
  INVX4 U496 ( .A(n552), .Y(n555) );
  AND2X4 U497 ( .A(A[12]), .B(B[12]), .Y(n552) );
  INVX4 U498 ( .A(n553), .Y(n554) );
  OR2X4 U499 ( .A(n558), .B(n559), .Y(n553) );
  AND2X4 U500 ( .A(n560), .B(n561), .Y(n558) );
  OR2X4 U501 ( .A(n562), .B(n563), .Y(n452) );
  AND2X4 U502 ( .A(n564), .B(n565), .Y(n563) );
  AND2X4 U503 ( .A(n566), .B(n468), .Y(n565) );
  OR2X4 U504 ( .A(n567), .B(n568), .Y(n468) );
  OR2X4 U505 ( .A(n569), .B(n570), .Y(n566) );
  INVX4 U506 ( .A(n467), .Y(n564) );
  AND2X4 U507 ( .A(n467), .B(n571), .Y(n562) );
  OR2X4 U508 ( .A(n572), .B(n466), .Y(n571) );
  AND2X4 U509 ( .A(n568), .B(n567), .Y(n466) );
  AND2X4 U510 ( .A(n569), .B(n570), .Y(n572) );
  INVX4 U511 ( .A(n567), .Y(n570) );
  AND2X4 U512 ( .A(A[11]), .B(B[13]), .Y(n567) );
  INVX4 U513 ( .A(n568), .Y(n569) );
  OR2X4 U514 ( .A(n573), .B(n574), .Y(n568) );
  AND2X4 U515 ( .A(n575), .B(n576), .Y(n573) );
  OR2X4 U516 ( .A(n577), .B(n578), .Y(n467) );
  AND2X4 U517 ( .A(n579), .B(n580), .Y(n578) );
  OR2X4 U518 ( .A(n581), .B(n582), .Y(n580) );
  AND2X4 U519 ( .A(A[9]), .B(n583), .Y(n582) );
  OR2X4 U520 ( .A(n584), .B(n297), .Y(n583) );
  AND2X4 U521 ( .A(B[15]), .B(n477), .Y(n584) );
  AND2X4 U522 ( .A(A[10]), .B(n585), .Y(n581) );
  OR2X4 U523 ( .A(n586), .B(n293), .Y(n585) );
  AND2X4 U524 ( .A(B[14]), .B(n587), .Y(n586) );
  INVX4 U525 ( .A(n484), .Y(n579) );
  AND2X4 U526 ( .A(n588), .B(n484), .Y(n577) );
  OR2X4 U527 ( .A(n589), .B(n590), .Y(n484) );
  AND2X4 U528 ( .A(n591), .B(n592), .Y(n589) );
  OR2X4 U529 ( .A(A[8]), .B(A[9]), .Y(n591) );
  OR2X4 U530 ( .A(n482), .B(n593), .Y(n588) );
  AND2X4 U531 ( .A(n477), .B(n587), .Y(n593) );
  INVX4 U532 ( .A(A[10]), .Y(n477) );
  AND2X4 U533 ( .A(n594), .B(A[10]), .Y(n482) );
  AND2X4 U534 ( .A(n306), .B(A[9]), .Y(n594) );
  NOR2X4 U535 ( .A(n595), .B(n596), .Y(n500) );
  OR2X4 U536 ( .A(n597), .B(n598), .Y(n596) );
  AND2X4 U537 ( .A(n599), .B(n600), .Y(n595) );
  OR2X4 U538 ( .A(n494), .B(n496), .Y(n498) );
  AND2X4 U539 ( .A(n601), .B(n602), .Y(n399) );
  AND2X4 U540 ( .A(n603), .B(n602), .Y(Y[23]) );
  OR2X4 U541 ( .A(n604), .B(n605), .Y(n602) );
  AND2X4 U542 ( .A(n606), .B(n607), .Y(n604) );
  OR2X4 U543 ( .A(n608), .B(n609), .Y(n606) );
  OR2X4 U544 ( .A(n610), .B(n611), .Y(n603) );
  OR2X4 U545 ( .A(n612), .B(n613), .Y(n611) );
  AND2X4 U546 ( .A(n614), .B(n601), .Y(n613) );
  NAND2X4 U547 ( .A(n615), .B(n616), .Y(n601) );
  OR2X4 U548 ( .A(n616), .B(n615), .Y(n614) );
  INVX4 U549 ( .A(n605), .Y(n615) );
  OR2X4 U550 ( .A(n617), .B(n618), .Y(n605) );
  NOR2X4 U551 ( .A(n494), .B(n496), .Y(n618) );
  AND2X4 U552 ( .A(n496), .B(n494), .Y(n617) );
  OR2X4 U553 ( .A(n619), .B(n620), .Y(n494) );
  OR2X4 U554 ( .A(n621), .B(n622), .Y(n620) );
  AND2X4 U555 ( .A(n623), .B(n624), .Y(n622) );
  OR2X4 U556 ( .A(n625), .B(n597), .Y(n624) );
  NOR2X4 U557 ( .A(n626), .B(n627), .Y(n597) );
  AND2X4 U558 ( .A(n626), .B(n627), .Y(n625) );
  AND2X4 U559 ( .A(n628), .B(n599), .Y(n621) );
  AND2X4 U560 ( .A(n627), .B(n600), .Y(n628) );
  AND2X4 U561 ( .A(n598), .B(n626), .Y(n619) );
  INVX4 U562 ( .A(n600), .Y(n626) );
  OR2X4 U563 ( .A(n629), .B(n630), .Y(n600) );
  AND2X4 U564 ( .A(n631), .B(n632), .Y(n629) );
  NOR2X4 U565 ( .A(n623), .B(n627), .Y(n598) );
  OR2X4 U566 ( .A(n633), .B(n175), .Y(n627) );
  INVX4 U567 ( .A(n599), .Y(n623) );
  OR2X4 U568 ( .A(n634), .B(n635), .Y(n599) );
  AND2X4 U569 ( .A(n636), .B(n637), .Y(n635) );
  AND2X4 U570 ( .A(n638), .B(n516), .Y(n637) );
  OR2X4 U571 ( .A(n639), .B(n640), .Y(n516) );
  OR2X4 U572 ( .A(n641), .B(n642), .Y(n638) );
  INVX4 U573 ( .A(n515), .Y(n636) );
  AND2X4 U574 ( .A(n515), .B(n643), .Y(n634) );
  OR2X4 U575 ( .A(n644), .B(n514), .Y(n643) );
  AND2X4 U576 ( .A(n640), .B(n639), .Y(n514) );
  AND2X4 U577 ( .A(n641), .B(n642), .Y(n644) );
  INVX4 U578 ( .A(n639), .Y(n642) );
  AND2X4 U579 ( .A(B[9]), .B(A[14]), .Y(n639) );
  INVX4 U580 ( .A(n640), .Y(n641) );
  OR2X4 U581 ( .A(n645), .B(n646), .Y(n640) );
  AND2X4 U582 ( .A(n647), .B(n648), .Y(n645) );
  OR2X4 U583 ( .A(n649), .B(n650), .Y(n515) );
  AND2X4 U584 ( .A(n651), .B(n652), .Y(n650) );
  AND2X4 U585 ( .A(n653), .B(n531), .Y(n652) );
  OR2X4 U586 ( .A(n654), .B(n655), .Y(n531) );
  OR2X4 U587 ( .A(n656), .B(n657), .Y(n653) );
  INVX4 U588 ( .A(n530), .Y(n651) );
  AND2X4 U589 ( .A(n530), .B(n658), .Y(n649) );
  OR2X4 U590 ( .A(n659), .B(n529), .Y(n658) );
  AND2X4 U591 ( .A(n655), .B(n654), .Y(n529) );
  AND2X4 U592 ( .A(n656), .B(n657), .Y(n659) );
  INVX4 U593 ( .A(n654), .Y(n657) );
  AND2X4 U594 ( .A(A[13]), .B(B[10]), .Y(n654) );
  INVX4 U595 ( .A(n655), .Y(n656) );
  OR2X4 U596 ( .A(n660), .B(n661), .Y(n655) );
  AND2X4 U597 ( .A(n662), .B(n663), .Y(n660) );
  OR2X4 U598 ( .A(n664), .B(n665), .Y(n530) );
  AND2X4 U599 ( .A(n666), .B(n667), .Y(n665) );
  AND2X4 U600 ( .A(n668), .B(n546), .Y(n667) );
  OR2X4 U601 ( .A(n669), .B(n670), .Y(n546) );
  OR2X4 U602 ( .A(n671), .B(n672), .Y(n668) );
  INVX4 U603 ( .A(n545), .Y(n666) );
  AND2X4 U604 ( .A(n545), .B(n673), .Y(n664) );
  OR2X4 U605 ( .A(n674), .B(n544), .Y(n673) );
  AND2X4 U606 ( .A(n670), .B(n669), .Y(n544) );
  AND2X4 U607 ( .A(n671), .B(n672), .Y(n674) );
  INVX4 U608 ( .A(n669), .Y(n672) );
  AND2X4 U609 ( .A(A[12]), .B(B[11]), .Y(n669) );
  INVX4 U610 ( .A(n670), .Y(n671) );
  OR2X4 U611 ( .A(n675), .B(n676), .Y(n670) );
  AND2X4 U612 ( .A(n677), .B(n678), .Y(n675) );
  OR2X4 U613 ( .A(n679), .B(n680), .Y(n545) );
  AND2X4 U614 ( .A(n681), .B(n682), .Y(n680) );
  AND2X4 U615 ( .A(n683), .B(n561), .Y(n682) );
  OR2X4 U616 ( .A(n684), .B(n685), .Y(n561) );
  OR2X4 U617 ( .A(n686), .B(n687), .Y(n683) );
  INVX4 U618 ( .A(n560), .Y(n681) );
  AND2X4 U619 ( .A(n560), .B(n688), .Y(n679) );
  OR2X4 U620 ( .A(n689), .B(n559), .Y(n688) );
  AND2X4 U621 ( .A(n685), .B(n684), .Y(n559) );
  AND2X4 U622 ( .A(n686), .B(n687), .Y(n689) );
  INVX4 U623 ( .A(n684), .Y(n687) );
  AND2X4 U624 ( .A(A[11]), .B(B[12]), .Y(n684) );
  INVX4 U625 ( .A(n685), .Y(n686) );
  OR2X4 U626 ( .A(n690), .B(n691), .Y(n685) );
  AND2X4 U627 ( .A(n692), .B(n693), .Y(n690) );
  OR2X4 U628 ( .A(n694), .B(n695), .Y(n560) );
  AND2X4 U629 ( .A(n696), .B(n697), .Y(n695) );
  AND2X4 U630 ( .A(n698), .B(n576), .Y(n697) );
  OR2X4 U631 ( .A(n699), .B(n700), .Y(n576) );
  OR2X4 U632 ( .A(n701), .B(n702), .Y(n698) );
  INVX4 U633 ( .A(n575), .Y(n696) );
  AND2X4 U634 ( .A(n575), .B(n703), .Y(n694) );
  OR2X4 U635 ( .A(n704), .B(n574), .Y(n703) );
  AND2X4 U636 ( .A(n700), .B(n699), .Y(n574) );
  AND2X4 U637 ( .A(n701), .B(n702), .Y(n704) );
  INVX4 U638 ( .A(n699), .Y(n702) );
  AND2X4 U639 ( .A(A[10]), .B(B[13]), .Y(n699) );
  INVX4 U640 ( .A(n700), .Y(n701) );
  OR2X4 U641 ( .A(n705), .B(n706), .Y(n700) );
  AND2X4 U642 ( .A(n707), .B(n708), .Y(n705) );
  OR2X4 U643 ( .A(n709), .B(n710), .Y(n575) );
  AND2X4 U644 ( .A(n711), .B(n712), .Y(n710) );
  OR2X4 U645 ( .A(n713), .B(n714), .Y(n712) );
  AND2X4 U646 ( .A(A[9]), .B(n715), .Y(n714) );
  OR2X4 U647 ( .A(n716), .B(n293), .Y(n715) );
  AND2X4 U648 ( .A(B[14]), .B(n717), .Y(n716) );
  AND2X4 U649 ( .A(A[8]), .B(n718), .Y(n713) );
  OR2X4 U650 ( .A(n719), .B(n297), .Y(n718) );
  AND2X4 U651 ( .A(B[15]), .B(n587), .Y(n719) );
  INVX4 U652 ( .A(n592), .Y(n711) );
  AND2X4 U653 ( .A(n720), .B(n592), .Y(n709) );
  OR2X4 U654 ( .A(n721), .B(n722), .Y(n592) );
  AND2X4 U655 ( .A(n723), .B(n724), .Y(n721) );
  OR2X4 U656 ( .A(A[7]), .B(A[8]), .Y(n723) );
  OR2X4 U657 ( .A(n590), .B(n725), .Y(n720) );
  AND2X4 U658 ( .A(n717), .B(n587), .Y(n725) );
  INVX4 U659 ( .A(A[9]), .Y(n587) );
  AND2X4 U660 ( .A(n726), .B(n306), .Y(n590) );
  AND2X4 U661 ( .A(A[9]), .B(A[8]), .Y(n726) );
  NOR2X4 U662 ( .A(n727), .B(n728), .Y(n496) );
  AND2X4 U663 ( .A(n729), .B(n730), .Y(n727) );
  NOR2X4 U664 ( .A(n608), .B(n609), .Y(n610) );
  AND2X4 U665 ( .A(n731), .B(n732), .Y(Y[22]) );
  NAND2X4 U666 ( .A(n733), .B(n609), .Y(n732) );
  OR2X4 U667 ( .A(n609), .B(n733), .Y(n731) );
  OR2X4 U668 ( .A(n608), .B(n612), .Y(n733) );
  INVX4 U669 ( .A(n607), .Y(n612) );
  OR2X4 U670 ( .A(n734), .B(n735), .Y(n607) );
  OR2X4 U671 ( .A(n736), .B(n737), .Y(n735) );
  AND2X4 U672 ( .A(n738), .B(n737), .Y(n608) );
  OR2X4 U673 ( .A(n739), .B(n616), .Y(n737) );
  NOR2X4 U674 ( .A(n740), .B(n741), .Y(n616) );
  AND2X4 U675 ( .A(n740), .B(n741), .Y(n739) );
  NOR2X4 U676 ( .A(n742), .B(n743), .Y(n741) );
  AND2X4 U677 ( .A(n744), .B(n745), .Y(n743) );
  AND2X4 U678 ( .A(n746), .B(n730), .Y(n745) );
  OR2X4 U679 ( .A(n747), .B(n748), .Y(n730) );
  OR2X4 U680 ( .A(n749), .B(n750), .Y(n746) );
  INVX4 U681 ( .A(n729), .Y(n744) );
  AND2X4 U682 ( .A(n729), .B(n751), .Y(n742) );
  OR2X4 U683 ( .A(n752), .B(n728), .Y(n751) );
  AND2X4 U684 ( .A(n748), .B(n747), .Y(n728) );
  AND2X4 U685 ( .A(n749), .B(n750), .Y(n752) );
  INVX4 U686 ( .A(n747), .Y(n750) );
  AND2X4 U687 ( .A(B[7]), .B(A[15]), .Y(n747) );
  INVX4 U688 ( .A(n748), .Y(n749) );
  OR2X4 U689 ( .A(n753), .B(n754), .Y(n748) );
  AND2X4 U690 ( .A(n755), .B(n756), .Y(n753) );
  OR2X4 U691 ( .A(n757), .B(n758), .Y(n729) );
  AND2X4 U692 ( .A(n759), .B(n760), .Y(n758) );
  AND2X4 U693 ( .A(n761), .B(n632), .Y(n760) );
  OR2X4 U694 ( .A(n762), .B(n763), .Y(n632) );
  OR2X4 U695 ( .A(n764), .B(n765), .Y(n761) );
  INVX4 U696 ( .A(n631), .Y(n759) );
  AND2X4 U697 ( .A(n631), .B(n766), .Y(n757) );
  OR2X4 U698 ( .A(n767), .B(n630), .Y(n766) );
  AND2X4 U699 ( .A(n763), .B(n762), .Y(n630) );
  AND2X4 U700 ( .A(n764), .B(n765), .Y(n767) );
  INVX4 U701 ( .A(n762), .Y(n765) );
  AND2X4 U702 ( .A(B[8]), .B(A[14]), .Y(n762) );
  INVX4 U703 ( .A(n763), .Y(n764) );
  OR2X4 U704 ( .A(n768), .B(n769), .Y(n763) );
  AND2X4 U705 ( .A(n770), .B(n771), .Y(n768) );
  OR2X4 U706 ( .A(n772), .B(n773), .Y(n631) );
  AND2X4 U707 ( .A(n774), .B(n775), .Y(n773) );
  AND2X4 U708 ( .A(n776), .B(n648), .Y(n775) );
  OR2X4 U709 ( .A(n777), .B(n778), .Y(n648) );
  OR2X4 U710 ( .A(n779), .B(n780), .Y(n776) );
  INVX4 U711 ( .A(n647), .Y(n774) );
  AND2X4 U712 ( .A(n647), .B(n781), .Y(n772) );
  OR2X4 U713 ( .A(n782), .B(n646), .Y(n781) );
  AND2X4 U714 ( .A(n778), .B(n777), .Y(n646) );
  AND2X4 U715 ( .A(n779), .B(n780), .Y(n782) );
  INVX4 U716 ( .A(n777), .Y(n780) );
  AND2X4 U717 ( .A(B[9]), .B(A[13]), .Y(n777) );
  INVX4 U718 ( .A(n778), .Y(n779) );
  OR2X4 U719 ( .A(n783), .B(n784), .Y(n778) );
  AND2X4 U720 ( .A(n785), .B(n786), .Y(n783) );
  OR2X4 U721 ( .A(n787), .B(n788), .Y(n647) );
  AND2X4 U722 ( .A(n789), .B(n790), .Y(n788) );
  AND2X4 U723 ( .A(n791), .B(n663), .Y(n790) );
  OR2X4 U724 ( .A(n792), .B(n793), .Y(n663) );
  OR2X4 U725 ( .A(n794), .B(n795), .Y(n791) );
  INVX4 U726 ( .A(n662), .Y(n789) );
  AND2X4 U727 ( .A(n662), .B(n796), .Y(n787) );
  OR2X4 U728 ( .A(n797), .B(n661), .Y(n796) );
  AND2X4 U729 ( .A(n793), .B(n792), .Y(n661) );
  AND2X4 U730 ( .A(n794), .B(n795), .Y(n797) );
  INVX4 U731 ( .A(n792), .Y(n795) );
  AND2X4 U732 ( .A(A[12]), .B(B[10]), .Y(n792) );
  INVX4 U733 ( .A(n793), .Y(n794) );
  OR2X4 U734 ( .A(n798), .B(n799), .Y(n793) );
  AND2X4 U735 ( .A(n800), .B(n801), .Y(n798) );
  OR2X4 U736 ( .A(n802), .B(n803), .Y(n662) );
  AND2X4 U737 ( .A(n804), .B(n805), .Y(n803) );
  AND2X4 U738 ( .A(n806), .B(n678), .Y(n805) );
  OR2X4 U739 ( .A(n807), .B(n808), .Y(n678) );
  OR2X4 U740 ( .A(n809), .B(n810), .Y(n806) );
  INVX4 U741 ( .A(n677), .Y(n804) );
  AND2X4 U742 ( .A(n677), .B(n811), .Y(n802) );
  OR2X4 U743 ( .A(n812), .B(n676), .Y(n811) );
  AND2X4 U744 ( .A(n808), .B(n807), .Y(n676) );
  AND2X4 U745 ( .A(n809), .B(n810), .Y(n812) );
  INVX4 U746 ( .A(n807), .Y(n810) );
  AND2X4 U747 ( .A(A[11]), .B(B[11]), .Y(n807) );
  INVX4 U748 ( .A(n808), .Y(n809) );
  OR2X4 U749 ( .A(n813), .B(n814), .Y(n808) );
  AND2X4 U750 ( .A(n815), .B(n816), .Y(n813) );
  OR2X4 U751 ( .A(n817), .B(n818), .Y(n677) );
  AND2X4 U752 ( .A(n819), .B(n820), .Y(n818) );
  AND2X4 U753 ( .A(n821), .B(n693), .Y(n820) );
  OR2X4 U754 ( .A(n822), .B(n823), .Y(n693) );
  OR2X4 U755 ( .A(n824), .B(n825), .Y(n821) );
  INVX4 U756 ( .A(n692), .Y(n819) );
  AND2X4 U757 ( .A(n692), .B(n826), .Y(n817) );
  OR2X4 U758 ( .A(n827), .B(n691), .Y(n826) );
  AND2X4 U759 ( .A(n823), .B(n822), .Y(n691) );
  AND2X4 U760 ( .A(n824), .B(n825), .Y(n827) );
  INVX4 U761 ( .A(n822), .Y(n825) );
  AND2X4 U762 ( .A(A[10]), .B(B[12]), .Y(n822) );
  INVX4 U763 ( .A(n823), .Y(n824) );
  OR2X4 U764 ( .A(n828), .B(n829), .Y(n823) );
  AND2X4 U765 ( .A(n830), .B(n831), .Y(n828) );
  OR2X4 U766 ( .A(n832), .B(n833), .Y(n692) );
  AND2X4 U767 ( .A(n834), .B(n835), .Y(n833) );
  AND2X4 U768 ( .A(n836), .B(n708), .Y(n835) );
  OR2X4 U769 ( .A(n837), .B(n838), .Y(n708) );
  OR2X4 U770 ( .A(n839), .B(n840), .Y(n836) );
  INVX4 U771 ( .A(n707), .Y(n834) );
  AND2X4 U772 ( .A(n707), .B(n841), .Y(n832) );
  OR2X4 U773 ( .A(n842), .B(n706), .Y(n841) );
  AND2X4 U774 ( .A(n838), .B(n837), .Y(n706) );
  AND2X4 U775 ( .A(n839), .B(n840), .Y(n842) );
  INVX4 U776 ( .A(n837), .Y(n840) );
  AND2X4 U777 ( .A(A[9]), .B(B[13]), .Y(n837) );
  INVX4 U778 ( .A(n838), .Y(n839) );
  OR2X4 U779 ( .A(n843), .B(n844), .Y(n838) );
  AND2X4 U780 ( .A(n845), .B(n846), .Y(n843) );
  OR2X4 U781 ( .A(n847), .B(n848), .Y(n707) );
  AND2X4 U782 ( .A(n849), .B(n850), .Y(n848) );
  OR2X4 U783 ( .A(n851), .B(n852), .Y(n850) );
  AND2X4 U784 ( .A(A[8]), .B(n853), .Y(n852) );
  OR2X4 U785 ( .A(n854), .B(n293), .Y(n853) );
  AND2X4 U786 ( .A(B[14]), .B(n855), .Y(n854) );
  AND2X4 U787 ( .A(A[7]), .B(n856), .Y(n851) );
  OR2X4 U788 ( .A(n857), .B(n297), .Y(n856) );
  AND2X4 U789 ( .A(B[15]), .B(n717), .Y(n857) );
  INVX4 U790 ( .A(n724), .Y(n849) );
  AND2X4 U791 ( .A(n858), .B(n724), .Y(n847) );
  OR2X4 U792 ( .A(n859), .B(n860), .Y(n724) );
  AND2X4 U793 ( .A(n861), .B(n862), .Y(n859) );
  OR2X4 U794 ( .A(A[6]), .B(A[7]), .Y(n861) );
  OR2X4 U795 ( .A(n722), .B(n863), .Y(n858) );
  AND2X4 U796 ( .A(n855), .B(n717), .Y(n863) );
  INVX4 U797 ( .A(A[8]), .Y(n717) );
  AND2X4 U798 ( .A(n864), .B(n306), .Y(n722) );
  AND2X4 U799 ( .A(A[8]), .B(A[7]), .Y(n864) );
  NOR2X4 U800 ( .A(n865), .B(n866), .Y(n740) );
  OR2X4 U801 ( .A(n867), .B(n868), .Y(n866) );
  AND2X4 U802 ( .A(n869), .B(n870), .Y(n865) );
  OR2X4 U803 ( .A(n734), .B(n736), .Y(n738) );
  AND2X4 U804 ( .A(n871), .B(n872), .Y(n609) );
  AND2X4 U805 ( .A(n873), .B(n872), .Y(Y[21]) );
  OR2X4 U806 ( .A(n874), .B(n875), .Y(n872) );
  AND2X4 U807 ( .A(n876), .B(n877), .Y(n874) );
  OR2X4 U808 ( .A(n878), .B(n879), .Y(n876) );
  OR2X4 U809 ( .A(n880), .B(n881), .Y(n873) );
  OR2X4 U810 ( .A(n882), .B(n883), .Y(n881) );
  AND2X4 U811 ( .A(n884), .B(n871), .Y(n883) );
  NAND2X4 U812 ( .A(n885), .B(n886), .Y(n871) );
  OR2X4 U813 ( .A(n886), .B(n885), .Y(n884) );
  INVX4 U814 ( .A(n875), .Y(n885) );
  OR2X4 U815 ( .A(n887), .B(n888), .Y(n875) );
  NOR2X4 U816 ( .A(n734), .B(n736), .Y(n888) );
  AND2X4 U817 ( .A(n736), .B(n734), .Y(n887) );
  OR2X4 U818 ( .A(n889), .B(n890), .Y(n734) );
  OR2X4 U819 ( .A(n891), .B(n892), .Y(n890) );
  AND2X4 U820 ( .A(n893), .B(n894), .Y(n892) );
  OR2X4 U821 ( .A(n895), .B(n867), .Y(n894) );
  NOR2X4 U822 ( .A(n896), .B(n897), .Y(n867) );
  AND2X4 U823 ( .A(n896), .B(n897), .Y(n895) );
  AND2X4 U824 ( .A(n898), .B(n869), .Y(n891) );
  AND2X4 U825 ( .A(n897), .B(n870), .Y(n898) );
  AND2X4 U826 ( .A(n868), .B(n896), .Y(n889) );
  INVX4 U827 ( .A(n870), .Y(n896) );
  OR2X4 U828 ( .A(n899), .B(n900), .Y(n870) );
  AND2X4 U829 ( .A(n901), .B(n902), .Y(n899) );
  NOR2X4 U830 ( .A(n893), .B(n897), .Y(n868) );
  OR2X4 U831 ( .A(n903), .B(n175), .Y(n897) );
  INVX4 U832 ( .A(n869), .Y(n893) );
  OR2X4 U833 ( .A(n904), .B(n905), .Y(n869) );
  AND2X4 U834 ( .A(n906), .B(n907), .Y(n905) );
  AND2X4 U835 ( .A(n908), .B(n756), .Y(n907) );
  OR2X4 U836 ( .A(n909), .B(n910), .Y(n756) );
  OR2X4 U837 ( .A(n911), .B(n912), .Y(n908) );
  INVX4 U838 ( .A(n755), .Y(n906) );
  AND2X4 U839 ( .A(n755), .B(n913), .Y(n904) );
  OR2X4 U840 ( .A(n914), .B(n754), .Y(n913) );
  AND2X4 U841 ( .A(n910), .B(n909), .Y(n754) );
  AND2X4 U842 ( .A(n911), .B(n912), .Y(n914) );
  INVX4 U843 ( .A(n909), .Y(n912) );
  AND2X4 U844 ( .A(B[7]), .B(A[14]), .Y(n909) );
  INVX4 U845 ( .A(n910), .Y(n911) );
  OR2X4 U846 ( .A(n915), .B(n916), .Y(n910) );
  AND2X4 U847 ( .A(n917), .B(n918), .Y(n915) );
  OR2X4 U848 ( .A(n919), .B(n920), .Y(n755) );
  AND2X4 U849 ( .A(n921), .B(n922), .Y(n920) );
  AND2X4 U850 ( .A(n923), .B(n771), .Y(n922) );
  OR2X4 U851 ( .A(n924), .B(n925), .Y(n771) );
  OR2X4 U852 ( .A(n926), .B(n927), .Y(n923) );
  INVX4 U853 ( .A(n770), .Y(n921) );
  AND2X4 U854 ( .A(n770), .B(n928), .Y(n919) );
  OR2X4 U855 ( .A(n929), .B(n769), .Y(n928) );
  AND2X4 U856 ( .A(n925), .B(n924), .Y(n769) );
  AND2X4 U857 ( .A(n926), .B(n927), .Y(n929) );
  INVX4 U858 ( .A(n924), .Y(n927) );
  AND2X4 U859 ( .A(B[8]), .B(A[13]), .Y(n924) );
  INVX4 U860 ( .A(n925), .Y(n926) );
  OR2X4 U861 ( .A(n930), .B(n931), .Y(n925) );
  AND2X4 U862 ( .A(n932), .B(n933), .Y(n930) );
  OR2X4 U863 ( .A(n934), .B(n935), .Y(n770) );
  AND2X4 U864 ( .A(n936), .B(n937), .Y(n935) );
  AND2X4 U865 ( .A(n938), .B(n786), .Y(n937) );
  OR2X4 U866 ( .A(n939), .B(n940), .Y(n786) );
  OR2X4 U867 ( .A(n941), .B(n942), .Y(n938) );
  INVX4 U868 ( .A(n785), .Y(n936) );
  AND2X4 U869 ( .A(n785), .B(n943), .Y(n934) );
  OR2X4 U870 ( .A(n944), .B(n784), .Y(n943) );
  AND2X4 U871 ( .A(n940), .B(n939), .Y(n784) );
  AND2X4 U872 ( .A(n941), .B(n942), .Y(n944) );
  INVX4 U873 ( .A(n939), .Y(n942) );
  AND2X4 U874 ( .A(B[9]), .B(A[12]), .Y(n939) );
  INVX4 U875 ( .A(n940), .Y(n941) );
  OR2X4 U876 ( .A(n945), .B(n946), .Y(n940) );
  AND2X4 U877 ( .A(n947), .B(n948), .Y(n945) );
  OR2X4 U878 ( .A(n949), .B(n950), .Y(n785) );
  AND2X4 U879 ( .A(n951), .B(n952), .Y(n950) );
  AND2X4 U880 ( .A(n953), .B(n801), .Y(n952) );
  OR2X4 U881 ( .A(n954), .B(n955), .Y(n801) );
  OR2X4 U882 ( .A(n956), .B(n957), .Y(n953) );
  INVX4 U883 ( .A(n800), .Y(n951) );
  AND2X4 U884 ( .A(n800), .B(n958), .Y(n949) );
  OR2X4 U885 ( .A(n959), .B(n799), .Y(n958) );
  AND2X4 U886 ( .A(n955), .B(n954), .Y(n799) );
  AND2X4 U887 ( .A(n956), .B(n957), .Y(n959) );
  INVX4 U888 ( .A(n954), .Y(n957) );
  AND2X4 U889 ( .A(A[11]), .B(B[10]), .Y(n954) );
  INVX4 U890 ( .A(n955), .Y(n956) );
  OR2X4 U891 ( .A(n960), .B(n961), .Y(n955) );
  AND2X4 U892 ( .A(n962), .B(n963), .Y(n960) );
  OR2X4 U893 ( .A(n964), .B(n965), .Y(n800) );
  AND2X4 U894 ( .A(n966), .B(n967), .Y(n965) );
  AND2X4 U895 ( .A(n968), .B(n816), .Y(n967) );
  OR2X4 U896 ( .A(n969), .B(n970), .Y(n816) );
  OR2X4 U897 ( .A(n971), .B(n972), .Y(n968) );
  INVX4 U898 ( .A(n815), .Y(n966) );
  AND2X4 U899 ( .A(n815), .B(n973), .Y(n964) );
  OR2X4 U900 ( .A(n974), .B(n814), .Y(n973) );
  AND2X4 U901 ( .A(n970), .B(n969), .Y(n814) );
  AND2X4 U902 ( .A(n971), .B(n972), .Y(n974) );
  INVX4 U903 ( .A(n969), .Y(n972) );
  AND2X4 U904 ( .A(A[10]), .B(B[11]), .Y(n969) );
  INVX4 U905 ( .A(n970), .Y(n971) );
  OR2X4 U906 ( .A(n975), .B(n976), .Y(n970) );
  AND2X4 U907 ( .A(n977), .B(n978), .Y(n975) );
  OR2X4 U908 ( .A(n979), .B(n980), .Y(n815) );
  AND2X4 U909 ( .A(n981), .B(n982), .Y(n980) );
  AND2X4 U910 ( .A(n983), .B(n831), .Y(n982) );
  OR2X4 U911 ( .A(n984), .B(n985), .Y(n831) );
  OR2X4 U912 ( .A(n986), .B(n987), .Y(n983) );
  INVX4 U913 ( .A(n830), .Y(n981) );
  AND2X4 U914 ( .A(n830), .B(n988), .Y(n979) );
  OR2X4 U915 ( .A(n989), .B(n829), .Y(n988) );
  AND2X4 U916 ( .A(n985), .B(n984), .Y(n829) );
  AND2X4 U917 ( .A(n986), .B(n987), .Y(n989) );
  INVX4 U918 ( .A(n984), .Y(n987) );
  AND2X4 U919 ( .A(A[9]), .B(B[12]), .Y(n984) );
  INVX4 U920 ( .A(n985), .Y(n986) );
  OR2X4 U921 ( .A(n990), .B(n991), .Y(n985) );
  AND2X4 U922 ( .A(n992), .B(n993), .Y(n990) );
  OR2X4 U923 ( .A(n994), .B(n995), .Y(n830) );
  AND2X4 U924 ( .A(n996), .B(n997), .Y(n995) );
  AND2X4 U925 ( .A(n998), .B(n846), .Y(n997) );
  OR2X4 U926 ( .A(n999), .B(n1000), .Y(n846) );
  OR2X4 U927 ( .A(n1001), .B(n1002), .Y(n998) );
  INVX4 U928 ( .A(n845), .Y(n996) );
  AND2X4 U929 ( .A(n845), .B(n1003), .Y(n994) );
  OR2X4 U930 ( .A(n1004), .B(n844), .Y(n1003) );
  AND2X4 U931 ( .A(n1000), .B(n999), .Y(n844) );
  AND2X4 U932 ( .A(n1001), .B(n1002), .Y(n1004) );
  INVX4 U933 ( .A(n999), .Y(n1002) );
  AND2X4 U934 ( .A(A[8]), .B(B[13]), .Y(n999) );
  INVX4 U935 ( .A(n1000), .Y(n1001) );
  OR2X4 U936 ( .A(n1005), .B(n1006), .Y(n1000) );
  AND2X4 U937 ( .A(n1007), .B(n1008), .Y(n1005) );
  OR2X4 U938 ( .A(n1009), .B(n1010), .Y(n845) );
  AND2X4 U939 ( .A(n1011), .B(n1012), .Y(n1010) );
  OR2X4 U940 ( .A(n1013), .B(n1014), .Y(n1012) );
  AND2X4 U941 ( .A(A[7]), .B(n1015), .Y(n1014) );
  OR2X4 U942 ( .A(n1016), .B(n293), .Y(n1015) );
  AND2X4 U943 ( .A(B[14]), .B(n1017), .Y(n1016) );
  AND2X4 U944 ( .A(A[6]), .B(n1018), .Y(n1013) );
  OR2X4 U945 ( .A(n1019), .B(n297), .Y(n1018) );
  AND2X4 U946 ( .A(B[15]), .B(n855), .Y(n1019) );
  INVX4 U947 ( .A(n862), .Y(n1011) );
  AND2X4 U948 ( .A(n1020), .B(n862), .Y(n1009) );
  OR2X4 U949 ( .A(n1021), .B(n1022), .Y(n862) );
  AND2X4 U950 ( .A(n1023), .B(n1024), .Y(n1021) );
  OR2X4 U951 ( .A(A[5]), .B(A[6]), .Y(n1023) );
  OR2X4 U952 ( .A(n860), .B(n1025), .Y(n1020) );
  AND2X4 U953 ( .A(n1017), .B(n855), .Y(n1025) );
  INVX4 U954 ( .A(A[7]), .Y(n855) );
  AND2X4 U955 ( .A(n1026), .B(n306), .Y(n860) );
  AND2X4 U956 ( .A(A[7]), .B(A[6]), .Y(n1026) );
  NOR2X4 U957 ( .A(n1027), .B(n1028), .Y(n736) );
  AND2X4 U958 ( .A(n1029), .B(n1030), .Y(n1027) );
  NOR2X4 U959 ( .A(n878), .B(n879), .Y(n880) );
  AND2X4 U960 ( .A(n1031), .B(n1032), .Y(Y[20]) );
  NAND2X4 U961 ( .A(n1033), .B(n879), .Y(n1032) );
  OR2X4 U962 ( .A(n879), .B(n1033), .Y(n1031) );
  OR2X4 U963 ( .A(n878), .B(n882), .Y(n1033) );
  INVX4 U964 ( .A(n877), .Y(n882) );
  OR2X4 U965 ( .A(n1034), .B(n1035), .Y(n877) );
  OR2X4 U966 ( .A(n1036), .B(n1037), .Y(n1035) );
  AND2X4 U967 ( .A(n1038), .B(n1037), .Y(n878) );
  OR2X4 U968 ( .A(n1039), .B(n886), .Y(n1037) );
  NOR2X4 U969 ( .A(n1040), .B(n1041), .Y(n886) );
  AND2X4 U970 ( .A(n1040), .B(n1041), .Y(n1039) );
  NOR2X4 U971 ( .A(n1042), .B(n1043), .Y(n1041) );
  AND2X4 U972 ( .A(n1044), .B(n1045), .Y(n1043) );
  AND2X4 U973 ( .A(n1046), .B(n1030), .Y(n1045) );
  OR2X4 U974 ( .A(n1047), .B(n1048), .Y(n1030) );
  OR2X4 U975 ( .A(n1049), .B(n1050), .Y(n1046) );
  INVX4 U976 ( .A(n1029), .Y(n1044) );
  AND2X4 U977 ( .A(n1029), .B(n1051), .Y(n1042) );
  OR2X4 U978 ( .A(n1052), .B(n1028), .Y(n1051) );
  AND2X4 U979 ( .A(n1048), .B(n1047), .Y(n1028) );
  AND2X4 U980 ( .A(n1049), .B(n1050), .Y(n1052) );
  INVX4 U981 ( .A(n1047), .Y(n1050) );
  AND2X4 U982 ( .A(B[5]), .B(A[15]), .Y(n1047) );
  INVX4 U983 ( .A(n1048), .Y(n1049) );
  OR2X4 U984 ( .A(n1053), .B(n1054), .Y(n1048) );
  AND2X4 U985 ( .A(n1055), .B(n1056), .Y(n1053) );
  OR2X4 U986 ( .A(n1057), .B(n1058), .Y(n1029) );
  AND2X4 U987 ( .A(n1059), .B(n1060), .Y(n1058) );
  AND2X4 U988 ( .A(n1061), .B(n902), .Y(n1060) );
  OR2X4 U989 ( .A(n1062), .B(n1063), .Y(n902) );
  OR2X4 U990 ( .A(n1064), .B(n1065), .Y(n1061) );
  INVX4 U991 ( .A(n901), .Y(n1059) );
  AND2X4 U992 ( .A(n901), .B(n1066), .Y(n1057) );
  OR2X4 U993 ( .A(n1067), .B(n900), .Y(n1066) );
  AND2X4 U994 ( .A(n1063), .B(n1062), .Y(n900) );
  AND2X4 U995 ( .A(n1064), .B(n1065), .Y(n1067) );
  INVX4 U996 ( .A(n1062), .Y(n1065) );
  AND2X4 U997 ( .A(B[6]), .B(A[14]), .Y(n1062) );
  INVX4 U998 ( .A(n1063), .Y(n1064) );
  OR2X4 U999 ( .A(n1068), .B(n1069), .Y(n1063) );
  AND2X4 U1000 ( .A(n1070), .B(n1071), .Y(n1068) );
  OR2X4 U1001 ( .A(n1072), .B(n1073), .Y(n901) );
  AND2X4 U1002 ( .A(n1074), .B(n1075), .Y(n1073) );
  AND2X4 U1003 ( .A(n1076), .B(n918), .Y(n1075) );
  OR2X4 U1004 ( .A(n1077), .B(n1078), .Y(n918) );
  OR2X4 U1005 ( .A(n1079), .B(n1080), .Y(n1076) );
  INVX4 U1006 ( .A(n917), .Y(n1074) );
  AND2X4 U1007 ( .A(n917), .B(n1081), .Y(n1072) );
  OR2X4 U1008 ( .A(n1082), .B(n916), .Y(n1081) );
  AND2X4 U1009 ( .A(n1078), .B(n1077), .Y(n916) );
  AND2X4 U1010 ( .A(n1079), .B(n1080), .Y(n1082) );
  INVX4 U1011 ( .A(n1077), .Y(n1080) );
  AND2X4 U1012 ( .A(B[7]), .B(A[13]), .Y(n1077) );
  INVX4 U1013 ( .A(n1078), .Y(n1079) );
  OR2X4 U1014 ( .A(n1083), .B(n1084), .Y(n1078) );
  AND2X4 U1015 ( .A(n1085), .B(n1086), .Y(n1083) );
  OR2X4 U1016 ( .A(n1087), .B(n1088), .Y(n917) );
  AND2X4 U1017 ( .A(n1089), .B(n1090), .Y(n1088) );
  AND2X4 U1018 ( .A(n1091), .B(n933), .Y(n1090) );
  OR2X4 U1019 ( .A(n1092), .B(n1093), .Y(n933) );
  OR2X4 U1020 ( .A(n1094), .B(n1095), .Y(n1091) );
  INVX4 U1021 ( .A(n932), .Y(n1089) );
  AND2X4 U1022 ( .A(n932), .B(n1096), .Y(n1087) );
  OR2X4 U1023 ( .A(n1097), .B(n931), .Y(n1096) );
  AND2X4 U1024 ( .A(n1093), .B(n1092), .Y(n931) );
  AND2X4 U1025 ( .A(n1094), .B(n1095), .Y(n1097) );
  INVX4 U1026 ( .A(n1092), .Y(n1095) );
  AND2X4 U1027 ( .A(B[8]), .B(A[12]), .Y(n1092) );
  INVX4 U1028 ( .A(n1093), .Y(n1094) );
  OR2X4 U1029 ( .A(n1098), .B(n1099), .Y(n1093) );
  AND2X4 U1030 ( .A(n1100), .B(n1101), .Y(n1098) );
  OR2X4 U1031 ( .A(n1102), .B(n1103), .Y(n932) );
  AND2X4 U1032 ( .A(n1104), .B(n1105), .Y(n1103) );
  AND2X4 U1033 ( .A(n1106), .B(n948), .Y(n1105) );
  OR2X4 U1034 ( .A(n1107), .B(n1108), .Y(n948) );
  OR2X4 U1035 ( .A(n1109), .B(n1110), .Y(n1106) );
  INVX4 U1036 ( .A(n947), .Y(n1104) );
  AND2X4 U1037 ( .A(n947), .B(n1111), .Y(n1102) );
  OR2X4 U1038 ( .A(n1112), .B(n946), .Y(n1111) );
  AND2X4 U1039 ( .A(n1108), .B(n1107), .Y(n946) );
  AND2X4 U1040 ( .A(n1109), .B(n1110), .Y(n1112) );
  INVX4 U1041 ( .A(n1107), .Y(n1110) );
  AND2X4 U1042 ( .A(B[9]), .B(A[11]), .Y(n1107) );
  INVX4 U1043 ( .A(n1108), .Y(n1109) );
  OR2X4 U1044 ( .A(n1113), .B(n1114), .Y(n1108) );
  AND2X4 U1045 ( .A(n1115), .B(n1116), .Y(n1113) );
  OR2X4 U1046 ( .A(n1117), .B(n1118), .Y(n947) );
  AND2X4 U1047 ( .A(n1119), .B(n1120), .Y(n1118) );
  AND2X4 U1048 ( .A(n1121), .B(n963), .Y(n1120) );
  OR2X4 U1049 ( .A(n1122), .B(n1123), .Y(n963) );
  OR2X4 U1050 ( .A(n1124), .B(n1125), .Y(n1121) );
  INVX4 U1051 ( .A(n962), .Y(n1119) );
  AND2X4 U1052 ( .A(n962), .B(n1126), .Y(n1117) );
  OR2X4 U1053 ( .A(n1127), .B(n961), .Y(n1126) );
  AND2X4 U1054 ( .A(n1123), .B(n1122), .Y(n961) );
  AND2X4 U1055 ( .A(n1124), .B(n1125), .Y(n1127) );
  INVX4 U1056 ( .A(n1122), .Y(n1125) );
  AND2X4 U1057 ( .A(A[10]), .B(B[10]), .Y(n1122) );
  INVX4 U1058 ( .A(n1123), .Y(n1124) );
  OR2X4 U1059 ( .A(n1128), .B(n1129), .Y(n1123) );
  AND2X4 U1060 ( .A(n1130), .B(n1131), .Y(n1128) );
  OR2X4 U1061 ( .A(n1132), .B(n1133), .Y(n962) );
  AND2X4 U1062 ( .A(n1134), .B(n1135), .Y(n1133) );
  AND2X4 U1063 ( .A(n1136), .B(n978), .Y(n1135) );
  OR2X4 U1064 ( .A(n1137), .B(n1138), .Y(n978) );
  OR2X4 U1065 ( .A(n1139), .B(n1140), .Y(n1136) );
  INVX4 U1066 ( .A(n977), .Y(n1134) );
  AND2X4 U1067 ( .A(n977), .B(n1141), .Y(n1132) );
  OR2X4 U1068 ( .A(n1142), .B(n976), .Y(n1141) );
  AND2X4 U1069 ( .A(n1138), .B(n1137), .Y(n976) );
  AND2X4 U1070 ( .A(n1139), .B(n1140), .Y(n1142) );
  INVX4 U1071 ( .A(n1137), .Y(n1140) );
  AND2X4 U1072 ( .A(A[9]), .B(B[11]), .Y(n1137) );
  INVX4 U1073 ( .A(n1138), .Y(n1139) );
  OR2X4 U1074 ( .A(n1143), .B(n1144), .Y(n1138) );
  AND2X4 U1075 ( .A(n1145), .B(n1146), .Y(n1143) );
  OR2X4 U1076 ( .A(n1147), .B(n1148), .Y(n977) );
  AND2X4 U1077 ( .A(n1149), .B(n1150), .Y(n1148) );
  AND2X4 U1078 ( .A(n1151), .B(n993), .Y(n1150) );
  OR2X4 U1079 ( .A(n1152), .B(n1153), .Y(n993) );
  OR2X4 U1080 ( .A(n1154), .B(n1155), .Y(n1151) );
  INVX4 U1081 ( .A(n992), .Y(n1149) );
  AND2X4 U1082 ( .A(n992), .B(n1156), .Y(n1147) );
  OR2X4 U1083 ( .A(n1157), .B(n991), .Y(n1156) );
  AND2X4 U1084 ( .A(n1153), .B(n1152), .Y(n991) );
  AND2X4 U1085 ( .A(n1154), .B(n1155), .Y(n1157) );
  INVX4 U1086 ( .A(n1152), .Y(n1155) );
  AND2X4 U1087 ( .A(A[8]), .B(B[12]), .Y(n1152) );
  INVX4 U1088 ( .A(n1153), .Y(n1154) );
  OR2X4 U1089 ( .A(n1158), .B(n1159), .Y(n1153) );
  AND2X4 U1090 ( .A(n1160), .B(n1161), .Y(n1158) );
  OR2X4 U1091 ( .A(n1162), .B(n1163), .Y(n992) );
  AND2X4 U1092 ( .A(n1164), .B(n1165), .Y(n1163) );
  AND2X4 U1093 ( .A(n1166), .B(n1008), .Y(n1165) );
  OR2X4 U1094 ( .A(n1167), .B(n1168), .Y(n1008) );
  OR2X4 U1095 ( .A(n1169), .B(n1170), .Y(n1166) );
  INVX4 U1096 ( .A(n1007), .Y(n1164) );
  AND2X4 U1097 ( .A(n1007), .B(n1171), .Y(n1162) );
  OR2X4 U1098 ( .A(n1172), .B(n1006), .Y(n1171) );
  AND2X4 U1099 ( .A(n1168), .B(n1167), .Y(n1006) );
  AND2X4 U1100 ( .A(n1169), .B(n1170), .Y(n1172) );
  INVX4 U1101 ( .A(n1167), .Y(n1170) );
  AND2X4 U1102 ( .A(A[7]), .B(B[13]), .Y(n1167) );
  INVX4 U1103 ( .A(n1168), .Y(n1169) );
  OR2X4 U1104 ( .A(n1173), .B(n1174), .Y(n1168) );
  AND2X4 U1105 ( .A(n1175), .B(n1176), .Y(n1173) );
  OR2X4 U1106 ( .A(n1177), .B(n1178), .Y(n1007) );
  AND2X4 U1107 ( .A(n1179), .B(n1180), .Y(n1178) );
  OR2X4 U1108 ( .A(n1181), .B(n1182), .Y(n1180) );
  AND2X4 U1109 ( .A(A[6]), .B(n1183), .Y(n1182) );
  OR2X4 U1110 ( .A(n1184), .B(n293), .Y(n1183) );
  AND2X4 U1111 ( .A(B[14]), .B(n1185), .Y(n1184) );
  AND2X4 U1112 ( .A(A[5]), .B(n1186), .Y(n1181) );
  OR2X4 U1113 ( .A(n1187), .B(n297), .Y(n1186) );
  AND2X4 U1114 ( .A(B[15]), .B(n1017), .Y(n1187) );
  INVX4 U1115 ( .A(n1024), .Y(n1179) );
  AND2X4 U1116 ( .A(n1188), .B(n1024), .Y(n1177) );
  OR2X4 U1117 ( .A(n1189), .B(n1190), .Y(n1024) );
  AND2X4 U1118 ( .A(n1191), .B(n1192), .Y(n1189) );
  OR2X4 U1119 ( .A(A[4]), .B(A[5]), .Y(n1191) );
  OR2X4 U1120 ( .A(n1022), .B(n1193), .Y(n1188) );
  AND2X4 U1121 ( .A(n1185), .B(n1017), .Y(n1193) );
  INVX4 U1122 ( .A(A[6]), .Y(n1017) );
  AND2X4 U1123 ( .A(n1194), .B(n306), .Y(n1022) );
  AND2X4 U1124 ( .A(A[6]), .B(A[5]), .Y(n1194) );
  NOR2X4 U1125 ( .A(n1195), .B(n1196), .Y(n1040) );
  OR2X4 U1126 ( .A(n1197), .B(n1198), .Y(n1196) );
  AND2X4 U1127 ( .A(n1199), .B(n1200), .Y(n1195) );
  OR2X4 U1128 ( .A(n1034), .B(n1036), .Y(n1038) );
  AND2X4 U1129 ( .A(n1201), .B(n1202), .Y(n879) );
  OR2X4 U1130 ( .A(n1203), .B(n1204), .Y(Y[1]) );
  AND2X4 U1131 ( .A(B[1]), .B(n1205), .Y(n1204) );
  OR2X4 U1132 ( .A(n1206), .B(n1207), .Y(n1205) );
  AND2X4 U1133 ( .A(A[0]), .B(n138), .Y(n1206) );
  INVX4 U1134 ( .A(B[0]), .Y(n138) );
  AND2X4 U1135 ( .A(B[0]), .B(n1208), .Y(n1203) );
  OR2X4 U1136 ( .A(n1209), .B(n1210), .Y(n1208) );
  AND2X4 U1137 ( .A(A[1]), .B(n132), .Y(n1209) );
  AND2X4 U1138 ( .A(n1211), .B(n1202), .Y(Y[19]) );
  OR2X4 U1139 ( .A(n1212), .B(n1213), .Y(n1202) );
  AND2X4 U1140 ( .A(n1214), .B(n1215), .Y(n1212) );
  OR2X4 U1141 ( .A(n1216), .B(n1217), .Y(n1214) );
  OR2X4 U1142 ( .A(n1218), .B(n1219), .Y(n1211) );
  OR2X4 U1143 ( .A(n1220), .B(n1221), .Y(n1219) );
  AND2X4 U1144 ( .A(n1222), .B(n1201), .Y(n1221) );
  NAND2X4 U1145 ( .A(n1223), .B(n1224), .Y(n1201) );
  OR2X4 U1146 ( .A(n1224), .B(n1223), .Y(n1222) );
  INVX4 U1147 ( .A(n1213), .Y(n1223) );
  OR2X4 U1148 ( .A(n1225), .B(n1226), .Y(n1213) );
  NOR2X4 U1149 ( .A(n1034), .B(n1036), .Y(n1226) );
  AND2X4 U1150 ( .A(n1036), .B(n1034), .Y(n1225) );
  OR2X4 U1151 ( .A(n1227), .B(n1228), .Y(n1034) );
  OR2X4 U1152 ( .A(n1229), .B(n1230), .Y(n1228) );
  AND2X4 U1153 ( .A(n1231), .B(n1232), .Y(n1230) );
  OR2X4 U1154 ( .A(n1233), .B(n1197), .Y(n1232) );
  NOR2X4 U1155 ( .A(n1234), .B(n1235), .Y(n1197) );
  AND2X4 U1156 ( .A(n1234), .B(n1235), .Y(n1233) );
  AND2X4 U1157 ( .A(n1236), .B(n1199), .Y(n1229) );
  AND2X4 U1158 ( .A(n1235), .B(n1200), .Y(n1236) );
  AND2X4 U1159 ( .A(n1198), .B(n1234), .Y(n1227) );
  INVX4 U1160 ( .A(n1200), .Y(n1234) );
  OR2X4 U1161 ( .A(n1237), .B(n1238), .Y(n1200) );
  AND2X4 U1162 ( .A(n1239), .B(n1240), .Y(n1237) );
  NOR2X4 U1163 ( .A(n1231), .B(n1235), .Y(n1198) );
  OR2X4 U1164 ( .A(n1241), .B(n175), .Y(n1235) );
  INVX4 U1165 ( .A(n1199), .Y(n1231) );
  OR2X4 U1166 ( .A(n1242), .B(n1243), .Y(n1199) );
  AND2X4 U1167 ( .A(n1244), .B(n1245), .Y(n1243) );
  AND2X4 U1168 ( .A(n1246), .B(n1056), .Y(n1245) );
  OR2X4 U1169 ( .A(n1247), .B(n1248), .Y(n1056) );
  OR2X4 U1170 ( .A(n1249), .B(n1250), .Y(n1246) );
  INVX4 U1171 ( .A(n1055), .Y(n1244) );
  AND2X4 U1172 ( .A(n1055), .B(n1251), .Y(n1242) );
  OR2X4 U1173 ( .A(n1252), .B(n1054), .Y(n1251) );
  AND2X4 U1174 ( .A(n1248), .B(n1247), .Y(n1054) );
  AND2X4 U1175 ( .A(n1249), .B(n1250), .Y(n1252) );
  INVX4 U1176 ( .A(n1247), .Y(n1250) );
  AND2X4 U1177 ( .A(B[5]), .B(A[14]), .Y(n1247) );
  INVX4 U1178 ( .A(n1248), .Y(n1249) );
  OR2X4 U1179 ( .A(n1253), .B(n1254), .Y(n1248) );
  AND2X4 U1180 ( .A(n1255), .B(n1256), .Y(n1253) );
  OR2X4 U1181 ( .A(n1257), .B(n1258), .Y(n1055) );
  AND2X4 U1182 ( .A(n1259), .B(n1260), .Y(n1258) );
  AND2X4 U1183 ( .A(n1261), .B(n1071), .Y(n1260) );
  OR2X4 U1184 ( .A(n1262), .B(n1263), .Y(n1071) );
  OR2X4 U1185 ( .A(n1264), .B(n1265), .Y(n1261) );
  INVX4 U1186 ( .A(n1070), .Y(n1259) );
  AND2X4 U1187 ( .A(n1070), .B(n1266), .Y(n1257) );
  OR2X4 U1188 ( .A(n1267), .B(n1069), .Y(n1266) );
  AND2X4 U1189 ( .A(n1263), .B(n1262), .Y(n1069) );
  AND2X4 U1190 ( .A(n1264), .B(n1265), .Y(n1267) );
  INVX4 U1191 ( .A(n1262), .Y(n1265) );
  AND2X4 U1192 ( .A(B[6]), .B(A[13]), .Y(n1262) );
  INVX4 U1193 ( .A(n1263), .Y(n1264) );
  OR2X4 U1194 ( .A(n1268), .B(n1269), .Y(n1263) );
  AND2X4 U1195 ( .A(n1270), .B(n1271), .Y(n1268) );
  OR2X4 U1196 ( .A(n1272), .B(n1273), .Y(n1070) );
  AND2X4 U1197 ( .A(n1274), .B(n1275), .Y(n1273) );
  AND2X4 U1198 ( .A(n1276), .B(n1086), .Y(n1275) );
  OR2X4 U1199 ( .A(n1277), .B(n1278), .Y(n1086) );
  OR2X4 U1200 ( .A(n1279), .B(n1280), .Y(n1276) );
  INVX4 U1201 ( .A(n1085), .Y(n1274) );
  AND2X4 U1202 ( .A(n1085), .B(n1281), .Y(n1272) );
  OR2X4 U1203 ( .A(n1282), .B(n1084), .Y(n1281) );
  AND2X4 U1204 ( .A(n1278), .B(n1277), .Y(n1084) );
  AND2X4 U1205 ( .A(n1279), .B(n1280), .Y(n1282) );
  INVX4 U1206 ( .A(n1277), .Y(n1280) );
  AND2X4 U1207 ( .A(B[7]), .B(A[12]), .Y(n1277) );
  INVX4 U1208 ( .A(n1278), .Y(n1279) );
  OR2X4 U1209 ( .A(n1283), .B(n1284), .Y(n1278) );
  AND2X4 U1210 ( .A(n1285), .B(n1286), .Y(n1283) );
  OR2X4 U1211 ( .A(n1287), .B(n1288), .Y(n1085) );
  AND2X4 U1212 ( .A(n1289), .B(n1290), .Y(n1288) );
  AND2X4 U1213 ( .A(n1291), .B(n1101), .Y(n1290) );
  OR2X4 U1214 ( .A(n1292), .B(n1293), .Y(n1101) );
  OR2X4 U1215 ( .A(n1294), .B(n1295), .Y(n1291) );
  INVX4 U1216 ( .A(n1100), .Y(n1289) );
  AND2X4 U1217 ( .A(n1100), .B(n1296), .Y(n1287) );
  OR2X4 U1218 ( .A(n1297), .B(n1099), .Y(n1296) );
  AND2X4 U1219 ( .A(n1293), .B(n1292), .Y(n1099) );
  AND2X4 U1220 ( .A(n1294), .B(n1295), .Y(n1297) );
  INVX4 U1221 ( .A(n1292), .Y(n1295) );
  AND2X4 U1222 ( .A(B[8]), .B(A[11]), .Y(n1292) );
  INVX4 U1223 ( .A(n1293), .Y(n1294) );
  OR2X4 U1224 ( .A(n1298), .B(n1299), .Y(n1293) );
  AND2X4 U1225 ( .A(n1300), .B(n1301), .Y(n1298) );
  OR2X4 U1226 ( .A(n1302), .B(n1303), .Y(n1100) );
  AND2X4 U1227 ( .A(n1304), .B(n1305), .Y(n1303) );
  AND2X4 U1228 ( .A(n1306), .B(n1116), .Y(n1305) );
  OR2X4 U1229 ( .A(n1307), .B(n1308), .Y(n1116) );
  OR2X4 U1230 ( .A(n1309), .B(n1310), .Y(n1306) );
  INVX4 U1231 ( .A(n1115), .Y(n1304) );
  AND2X4 U1232 ( .A(n1115), .B(n1311), .Y(n1302) );
  OR2X4 U1233 ( .A(n1312), .B(n1114), .Y(n1311) );
  AND2X4 U1234 ( .A(n1308), .B(n1307), .Y(n1114) );
  AND2X4 U1235 ( .A(n1309), .B(n1310), .Y(n1312) );
  INVX4 U1236 ( .A(n1307), .Y(n1310) );
  AND2X4 U1237 ( .A(B[9]), .B(A[10]), .Y(n1307) );
  INVX4 U1238 ( .A(n1308), .Y(n1309) );
  OR2X4 U1239 ( .A(n1313), .B(n1314), .Y(n1308) );
  AND2X4 U1240 ( .A(n1315), .B(n1316), .Y(n1313) );
  OR2X4 U1241 ( .A(n1317), .B(n1318), .Y(n1115) );
  AND2X4 U1242 ( .A(n1319), .B(n1320), .Y(n1318) );
  AND2X4 U1243 ( .A(n1321), .B(n1131), .Y(n1320) );
  OR2X4 U1244 ( .A(n1322), .B(n1323), .Y(n1131) );
  OR2X4 U1245 ( .A(n1324), .B(n1325), .Y(n1321) );
  INVX4 U1246 ( .A(n1130), .Y(n1319) );
  AND2X4 U1247 ( .A(n1130), .B(n1326), .Y(n1317) );
  OR2X4 U1248 ( .A(n1327), .B(n1129), .Y(n1326) );
  AND2X4 U1249 ( .A(n1323), .B(n1322), .Y(n1129) );
  AND2X4 U1250 ( .A(n1324), .B(n1325), .Y(n1327) );
  INVX4 U1251 ( .A(n1322), .Y(n1325) );
  AND2X4 U1252 ( .A(A[9]), .B(B[10]), .Y(n1322) );
  INVX4 U1253 ( .A(n1323), .Y(n1324) );
  OR2X4 U1254 ( .A(n1328), .B(n1329), .Y(n1323) );
  AND2X4 U1255 ( .A(n1330), .B(n1331), .Y(n1328) );
  OR2X4 U1256 ( .A(n1332), .B(n1333), .Y(n1130) );
  AND2X4 U1257 ( .A(n1334), .B(n1335), .Y(n1333) );
  AND2X4 U1258 ( .A(n1336), .B(n1146), .Y(n1335) );
  OR2X4 U1259 ( .A(n1337), .B(n1338), .Y(n1146) );
  OR2X4 U1260 ( .A(n1339), .B(n1340), .Y(n1336) );
  INVX4 U1261 ( .A(n1145), .Y(n1334) );
  AND2X4 U1262 ( .A(n1145), .B(n1341), .Y(n1332) );
  OR2X4 U1263 ( .A(n1342), .B(n1144), .Y(n1341) );
  AND2X4 U1264 ( .A(n1338), .B(n1337), .Y(n1144) );
  AND2X4 U1265 ( .A(n1339), .B(n1340), .Y(n1342) );
  INVX4 U1266 ( .A(n1337), .Y(n1340) );
  AND2X4 U1267 ( .A(A[8]), .B(B[11]), .Y(n1337) );
  INVX4 U1268 ( .A(n1338), .Y(n1339) );
  OR2X4 U1269 ( .A(n1343), .B(n1344), .Y(n1338) );
  AND2X4 U1270 ( .A(n1345), .B(n1346), .Y(n1343) );
  OR2X4 U1271 ( .A(n1347), .B(n1348), .Y(n1145) );
  AND2X4 U1272 ( .A(n1349), .B(n1350), .Y(n1348) );
  AND2X4 U1273 ( .A(n1351), .B(n1161), .Y(n1350) );
  OR2X4 U1274 ( .A(n1352), .B(n1353), .Y(n1161) );
  OR2X4 U1275 ( .A(n1354), .B(n1355), .Y(n1351) );
  INVX4 U1276 ( .A(n1160), .Y(n1349) );
  AND2X4 U1277 ( .A(n1160), .B(n1356), .Y(n1347) );
  OR2X4 U1278 ( .A(n1357), .B(n1159), .Y(n1356) );
  AND2X4 U1279 ( .A(n1353), .B(n1352), .Y(n1159) );
  AND2X4 U1280 ( .A(n1354), .B(n1355), .Y(n1357) );
  INVX4 U1281 ( .A(n1352), .Y(n1355) );
  AND2X4 U1282 ( .A(A[7]), .B(B[12]), .Y(n1352) );
  INVX4 U1283 ( .A(n1353), .Y(n1354) );
  OR2X4 U1284 ( .A(n1358), .B(n1359), .Y(n1353) );
  AND2X4 U1285 ( .A(n1360), .B(n1361), .Y(n1358) );
  OR2X4 U1286 ( .A(n1362), .B(n1363), .Y(n1160) );
  AND2X4 U1287 ( .A(n1364), .B(n1365), .Y(n1363) );
  AND2X4 U1288 ( .A(n1366), .B(n1176), .Y(n1365) );
  OR2X4 U1289 ( .A(n1367), .B(n1368), .Y(n1176) );
  OR2X4 U1290 ( .A(n1369), .B(n1370), .Y(n1366) );
  INVX4 U1291 ( .A(n1175), .Y(n1364) );
  AND2X4 U1292 ( .A(n1175), .B(n1371), .Y(n1362) );
  OR2X4 U1293 ( .A(n1372), .B(n1174), .Y(n1371) );
  AND2X4 U1294 ( .A(n1368), .B(n1367), .Y(n1174) );
  AND2X4 U1295 ( .A(n1369), .B(n1370), .Y(n1372) );
  INVX4 U1296 ( .A(n1367), .Y(n1370) );
  AND2X4 U1297 ( .A(A[6]), .B(B[13]), .Y(n1367) );
  INVX4 U1298 ( .A(n1368), .Y(n1369) );
  OR2X4 U1299 ( .A(n1373), .B(n1374), .Y(n1368) );
  AND2X4 U1300 ( .A(n1375), .B(n1376), .Y(n1373) );
  OR2X4 U1301 ( .A(n1377), .B(n1378), .Y(n1175) );
  AND2X4 U1302 ( .A(n1379), .B(n1380), .Y(n1378) );
  OR2X4 U1303 ( .A(n1381), .B(n1382), .Y(n1380) );
  AND2X4 U1304 ( .A(A[5]), .B(n1383), .Y(n1382) );
  OR2X4 U1305 ( .A(n1384), .B(n293), .Y(n1383) );
  AND2X4 U1306 ( .A(B[14]), .B(n1385), .Y(n1384) );
  AND2X4 U1307 ( .A(A[4]), .B(n1386), .Y(n1381) );
  OR2X4 U1308 ( .A(n1387), .B(n297), .Y(n1386) );
  AND2X4 U1309 ( .A(B[15]), .B(n1185), .Y(n1387) );
  INVX4 U1310 ( .A(n1192), .Y(n1379) );
  AND2X4 U1311 ( .A(n1388), .B(n1192), .Y(n1377) );
  OR2X4 U1312 ( .A(n1389), .B(n1390), .Y(n1192) );
  AND2X4 U1313 ( .A(n1391), .B(n1392), .Y(n1389) );
  OR2X4 U1314 ( .A(A[3]), .B(A[4]), .Y(n1391) );
  OR2X4 U1315 ( .A(n1190), .B(n1393), .Y(n1388) );
  AND2X4 U1316 ( .A(n1385), .B(n1185), .Y(n1393) );
  INVX4 U1317 ( .A(A[5]), .Y(n1185) );
  AND2X4 U1318 ( .A(n1394), .B(n306), .Y(n1190) );
  AND2X4 U1319 ( .A(A[5]), .B(A[4]), .Y(n1394) );
  NOR2X4 U1320 ( .A(n1395), .B(n1396), .Y(n1036) );
  AND2X4 U1321 ( .A(n1397), .B(n1398), .Y(n1395) );
  NOR2X4 U1322 ( .A(n1217), .B(n1216), .Y(n1218) );
  OR2X4 U1323 ( .A(n1399), .B(n1400), .Y(Y[18]) );
  AND2X4 U1324 ( .A(n1401), .B(n1217), .Y(n1400) );
  NOR2X4 U1325 ( .A(n1217), .B(n1401), .Y(n1399) );
  NOR2X4 U1326 ( .A(n1216), .B(n1220), .Y(n1401) );
  INVX4 U1327 ( .A(n1215), .Y(n1220) );
  OR2X4 U1328 ( .A(n1402), .B(n1403), .Y(n1215) );
  OR2X4 U1329 ( .A(n1404), .B(n1405), .Y(n1403) );
  AND2X4 U1330 ( .A(n1406), .B(n1405), .Y(n1216) );
  OR2X4 U1331 ( .A(n1407), .B(n1224), .Y(n1405) );
  NOR2X4 U1332 ( .A(n1408), .B(n1409), .Y(n1224) );
  AND2X4 U1333 ( .A(n1408), .B(n1409), .Y(n1407) );
  NOR2X4 U1334 ( .A(n1410), .B(n1411), .Y(n1409) );
  AND2X4 U1335 ( .A(n1412), .B(n1413), .Y(n1411) );
  AND2X4 U1336 ( .A(n1414), .B(n1398), .Y(n1413) );
  OR2X4 U1337 ( .A(n1415), .B(n1416), .Y(n1398) );
  OR2X4 U1338 ( .A(n1417), .B(n1418), .Y(n1414) );
  INVX4 U1339 ( .A(n1397), .Y(n1412) );
  AND2X4 U1340 ( .A(n1397), .B(n1419), .Y(n1410) );
  OR2X4 U1341 ( .A(n1420), .B(n1396), .Y(n1419) );
  AND2X4 U1342 ( .A(n1416), .B(n1415), .Y(n1396) );
  AND2X4 U1343 ( .A(n1417), .B(n1418), .Y(n1420) );
  INVX4 U1344 ( .A(n1415), .Y(n1418) );
  AND2X4 U1345 ( .A(B[3]), .B(A[15]), .Y(n1415) );
  INVX4 U1346 ( .A(n1416), .Y(n1417) );
  OR2X4 U1347 ( .A(n1421), .B(n1422), .Y(n1416) );
  AND2X4 U1348 ( .A(n1423), .B(n1424), .Y(n1421) );
  OR2X4 U1349 ( .A(n1425), .B(n1426), .Y(n1397) );
  AND2X4 U1350 ( .A(n1427), .B(n1428), .Y(n1426) );
  AND2X4 U1351 ( .A(n1429), .B(n1240), .Y(n1428) );
  OR2X4 U1352 ( .A(n1430), .B(n1431), .Y(n1240) );
  OR2X4 U1353 ( .A(n1432), .B(n1433), .Y(n1429) );
  INVX4 U1354 ( .A(n1239), .Y(n1427) );
  AND2X4 U1355 ( .A(n1239), .B(n1434), .Y(n1425) );
  OR2X4 U1356 ( .A(n1435), .B(n1238), .Y(n1434) );
  AND2X4 U1357 ( .A(n1431), .B(n1430), .Y(n1238) );
  AND2X4 U1358 ( .A(n1432), .B(n1433), .Y(n1435) );
  INVX4 U1359 ( .A(n1430), .Y(n1433) );
  AND2X4 U1360 ( .A(B[4]), .B(A[14]), .Y(n1430) );
  INVX4 U1361 ( .A(n1431), .Y(n1432) );
  OR2X4 U1362 ( .A(n1436), .B(n1437), .Y(n1431) );
  AND2X4 U1363 ( .A(n1438), .B(n1439), .Y(n1436) );
  OR2X4 U1364 ( .A(n1440), .B(n1441), .Y(n1239) );
  AND2X4 U1365 ( .A(n1442), .B(n1443), .Y(n1441) );
  AND2X4 U1366 ( .A(n1444), .B(n1256), .Y(n1443) );
  OR2X4 U1367 ( .A(n1445), .B(n1446), .Y(n1256) );
  OR2X4 U1368 ( .A(n1447), .B(n1448), .Y(n1444) );
  INVX4 U1369 ( .A(n1255), .Y(n1442) );
  AND2X4 U1370 ( .A(n1255), .B(n1449), .Y(n1440) );
  OR2X4 U1371 ( .A(n1450), .B(n1254), .Y(n1449) );
  AND2X4 U1372 ( .A(n1446), .B(n1445), .Y(n1254) );
  AND2X4 U1373 ( .A(n1447), .B(n1448), .Y(n1450) );
  INVX4 U1374 ( .A(n1445), .Y(n1448) );
  AND2X4 U1375 ( .A(B[5]), .B(A[13]), .Y(n1445) );
  INVX4 U1376 ( .A(n1446), .Y(n1447) );
  OR2X4 U1377 ( .A(n1451), .B(n1452), .Y(n1446) );
  AND2X4 U1378 ( .A(n1453), .B(n1454), .Y(n1451) );
  OR2X4 U1379 ( .A(n1455), .B(n1456), .Y(n1255) );
  AND2X4 U1380 ( .A(n1457), .B(n1458), .Y(n1456) );
  AND2X4 U1381 ( .A(n1459), .B(n1271), .Y(n1458) );
  OR2X4 U1382 ( .A(n1460), .B(n1461), .Y(n1271) );
  OR2X4 U1383 ( .A(n1462), .B(n1463), .Y(n1459) );
  INVX4 U1384 ( .A(n1270), .Y(n1457) );
  AND2X4 U1385 ( .A(n1270), .B(n1464), .Y(n1455) );
  OR2X4 U1386 ( .A(n1465), .B(n1269), .Y(n1464) );
  AND2X4 U1387 ( .A(n1461), .B(n1460), .Y(n1269) );
  AND2X4 U1388 ( .A(n1462), .B(n1463), .Y(n1465) );
  INVX4 U1389 ( .A(n1460), .Y(n1463) );
  AND2X4 U1390 ( .A(B[6]), .B(A[12]), .Y(n1460) );
  INVX4 U1391 ( .A(n1461), .Y(n1462) );
  OR2X4 U1392 ( .A(n1466), .B(n1467), .Y(n1461) );
  AND2X4 U1393 ( .A(n1468), .B(n1469), .Y(n1466) );
  OR2X4 U1394 ( .A(n1470), .B(n1471), .Y(n1270) );
  AND2X4 U1395 ( .A(n1472), .B(n1473), .Y(n1471) );
  AND2X4 U1396 ( .A(n1474), .B(n1286), .Y(n1473) );
  OR2X4 U1397 ( .A(n1475), .B(n1476), .Y(n1286) );
  OR2X4 U1398 ( .A(n1477), .B(n1478), .Y(n1474) );
  INVX4 U1399 ( .A(n1285), .Y(n1472) );
  AND2X4 U1400 ( .A(n1285), .B(n1479), .Y(n1470) );
  OR2X4 U1401 ( .A(n1480), .B(n1284), .Y(n1479) );
  AND2X4 U1402 ( .A(n1476), .B(n1475), .Y(n1284) );
  AND2X4 U1403 ( .A(n1477), .B(n1478), .Y(n1480) );
  INVX4 U1404 ( .A(n1475), .Y(n1478) );
  AND2X4 U1405 ( .A(B[7]), .B(A[11]), .Y(n1475) );
  INVX4 U1406 ( .A(n1476), .Y(n1477) );
  OR2X4 U1407 ( .A(n1481), .B(n1482), .Y(n1476) );
  AND2X4 U1408 ( .A(n1483), .B(n1484), .Y(n1481) );
  OR2X4 U1409 ( .A(n1485), .B(n1486), .Y(n1285) );
  AND2X4 U1410 ( .A(n1487), .B(n1488), .Y(n1486) );
  AND2X4 U1411 ( .A(n1489), .B(n1301), .Y(n1488) );
  OR2X4 U1412 ( .A(n1490), .B(n1491), .Y(n1301) );
  OR2X4 U1413 ( .A(n1492), .B(n1493), .Y(n1489) );
  INVX4 U1414 ( .A(n1300), .Y(n1487) );
  AND2X4 U1415 ( .A(n1300), .B(n1494), .Y(n1485) );
  OR2X4 U1416 ( .A(n1495), .B(n1299), .Y(n1494) );
  AND2X4 U1417 ( .A(n1491), .B(n1490), .Y(n1299) );
  AND2X4 U1418 ( .A(n1492), .B(n1493), .Y(n1495) );
  INVX4 U1419 ( .A(n1490), .Y(n1493) );
  AND2X4 U1420 ( .A(B[8]), .B(A[10]), .Y(n1490) );
  INVX4 U1421 ( .A(n1491), .Y(n1492) );
  OR2X4 U1422 ( .A(n1496), .B(n1497), .Y(n1491) );
  AND2X4 U1423 ( .A(n1498), .B(n1499), .Y(n1496) );
  OR2X4 U1424 ( .A(n1500), .B(n1501), .Y(n1300) );
  AND2X4 U1425 ( .A(n1502), .B(n1503), .Y(n1501) );
  AND2X4 U1426 ( .A(n1504), .B(n1316), .Y(n1503) );
  OR2X4 U1427 ( .A(n1505), .B(n1506), .Y(n1316) );
  OR2X4 U1428 ( .A(n1507), .B(n1508), .Y(n1504) );
  INVX4 U1429 ( .A(n1315), .Y(n1502) );
  AND2X4 U1430 ( .A(n1315), .B(n1509), .Y(n1500) );
  OR2X4 U1431 ( .A(n1510), .B(n1314), .Y(n1509) );
  AND2X4 U1432 ( .A(n1506), .B(n1505), .Y(n1314) );
  AND2X4 U1433 ( .A(n1507), .B(n1508), .Y(n1510) );
  INVX4 U1434 ( .A(n1505), .Y(n1508) );
  AND2X4 U1435 ( .A(B[9]), .B(A[9]), .Y(n1505) );
  INVX4 U1436 ( .A(n1506), .Y(n1507) );
  OR2X4 U1437 ( .A(n1511), .B(n1512), .Y(n1506) );
  AND2X4 U1438 ( .A(n1513), .B(n1514), .Y(n1511) );
  OR2X4 U1439 ( .A(n1515), .B(n1516), .Y(n1315) );
  AND2X4 U1440 ( .A(n1517), .B(n1518), .Y(n1516) );
  AND2X4 U1441 ( .A(n1519), .B(n1331), .Y(n1518) );
  OR2X4 U1442 ( .A(n1520), .B(n1521), .Y(n1331) );
  OR2X4 U1443 ( .A(n1522), .B(n1523), .Y(n1519) );
  INVX4 U1444 ( .A(n1330), .Y(n1517) );
  AND2X4 U1445 ( .A(n1330), .B(n1524), .Y(n1515) );
  OR2X4 U1446 ( .A(n1525), .B(n1329), .Y(n1524) );
  AND2X4 U1447 ( .A(n1521), .B(n1520), .Y(n1329) );
  AND2X4 U1448 ( .A(n1522), .B(n1523), .Y(n1525) );
  INVX4 U1449 ( .A(n1520), .Y(n1523) );
  AND2X4 U1450 ( .A(A[8]), .B(B[10]), .Y(n1520) );
  INVX4 U1451 ( .A(n1521), .Y(n1522) );
  OR2X4 U1452 ( .A(n1526), .B(n1527), .Y(n1521) );
  AND2X4 U1453 ( .A(n1528), .B(n1529), .Y(n1526) );
  OR2X4 U1454 ( .A(n1530), .B(n1531), .Y(n1330) );
  AND2X4 U1455 ( .A(n1532), .B(n1533), .Y(n1531) );
  AND2X4 U1456 ( .A(n1534), .B(n1346), .Y(n1533) );
  OR2X4 U1457 ( .A(n1535), .B(n1536), .Y(n1346) );
  OR2X4 U1458 ( .A(n1537), .B(n1538), .Y(n1534) );
  INVX4 U1459 ( .A(n1345), .Y(n1532) );
  AND2X4 U1460 ( .A(n1345), .B(n1539), .Y(n1530) );
  OR2X4 U1461 ( .A(n1540), .B(n1344), .Y(n1539) );
  AND2X4 U1462 ( .A(n1536), .B(n1535), .Y(n1344) );
  AND2X4 U1463 ( .A(n1537), .B(n1538), .Y(n1540) );
  INVX4 U1464 ( .A(n1535), .Y(n1538) );
  AND2X4 U1465 ( .A(A[7]), .B(B[11]), .Y(n1535) );
  INVX4 U1466 ( .A(n1536), .Y(n1537) );
  OR2X4 U1467 ( .A(n1541), .B(n1542), .Y(n1536) );
  AND2X4 U1468 ( .A(n1543), .B(n1544), .Y(n1541) );
  OR2X4 U1469 ( .A(n1545), .B(n1546), .Y(n1345) );
  AND2X4 U1470 ( .A(n1547), .B(n1548), .Y(n1546) );
  AND2X4 U1471 ( .A(n1549), .B(n1361), .Y(n1548) );
  OR2X4 U1472 ( .A(n1550), .B(n1551), .Y(n1361) );
  OR2X4 U1473 ( .A(n1552), .B(n1553), .Y(n1549) );
  INVX4 U1474 ( .A(n1360), .Y(n1547) );
  AND2X4 U1475 ( .A(n1360), .B(n1554), .Y(n1545) );
  OR2X4 U1476 ( .A(n1555), .B(n1359), .Y(n1554) );
  AND2X4 U1477 ( .A(n1551), .B(n1550), .Y(n1359) );
  AND2X4 U1478 ( .A(n1552), .B(n1553), .Y(n1555) );
  INVX4 U1479 ( .A(n1550), .Y(n1553) );
  AND2X4 U1480 ( .A(A[6]), .B(B[12]), .Y(n1550) );
  INVX4 U1481 ( .A(n1551), .Y(n1552) );
  OR2X4 U1482 ( .A(n1556), .B(n1557), .Y(n1551) );
  AND2X4 U1483 ( .A(n1558), .B(n1559), .Y(n1556) );
  OR2X4 U1484 ( .A(n1560), .B(n1561), .Y(n1360) );
  AND2X4 U1485 ( .A(n1562), .B(n1563), .Y(n1561) );
  AND2X4 U1486 ( .A(n1564), .B(n1376), .Y(n1563) );
  OR2X4 U1487 ( .A(n1565), .B(n1566), .Y(n1376) );
  OR2X4 U1488 ( .A(n1567), .B(n1568), .Y(n1564) );
  INVX4 U1489 ( .A(n1375), .Y(n1562) );
  AND2X4 U1490 ( .A(n1375), .B(n1569), .Y(n1560) );
  OR2X4 U1491 ( .A(n1570), .B(n1374), .Y(n1569) );
  AND2X4 U1492 ( .A(n1566), .B(n1565), .Y(n1374) );
  AND2X4 U1493 ( .A(n1567), .B(n1568), .Y(n1570) );
  INVX4 U1494 ( .A(n1565), .Y(n1568) );
  AND2X4 U1495 ( .A(A[5]), .B(B[13]), .Y(n1565) );
  INVX4 U1496 ( .A(n1566), .Y(n1567) );
  OR2X4 U1497 ( .A(n1571), .B(n1572), .Y(n1566) );
  AND2X4 U1498 ( .A(n1573), .B(n1574), .Y(n1571) );
  OR2X4 U1499 ( .A(n1575), .B(n1576), .Y(n1375) );
  AND2X4 U1500 ( .A(n1577), .B(n1578), .Y(n1576) );
  OR2X4 U1501 ( .A(n1579), .B(n1580), .Y(n1578) );
  AND2X4 U1502 ( .A(A[4]), .B(n1581), .Y(n1580) );
  OR2X4 U1503 ( .A(n1582), .B(n293), .Y(n1581) );
  AND2X4 U1504 ( .A(B[14]), .B(n1583), .Y(n1582) );
  AND2X4 U1505 ( .A(A[3]), .B(n1584), .Y(n1579) );
  OR2X4 U1506 ( .A(n1585), .B(n297), .Y(n1584) );
  AND2X4 U1507 ( .A(B[15]), .B(n1385), .Y(n1585) );
  INVX4 U1508 ( .A(n1392), .Y(n1577) );
  AND2X4 U1509 ( .A(n1586), .B(n1392), .Y(n1575) );
  OR2X4 U1510 ( .A(n1587), .B(n1588), .Y(n1392) );
  AND2X4 U1511 ( .A(n1589), .B(n1590), .Y(n1587) );
  OR2X4 U1512 ( .A(A[2]), .B(A[3]), .Y(n1590) );
  OR2X4 U1513 ( .A(n1390), .B(n1591), .Y(n1586) );
  AND2X4 U1514 ( .A(n1583), .B(n1385), .Y(n1591) );
  INVX4 U1515 ( .A(A[4]), .Y(n1385) );
  AND2X4 U1516 ( .A(n1592), .B(n306), .Y(n1390) );
  AND2X4 U1517 ( .A(A[4]), .B(A[3]), .Y(n1592) );
  NOR2X4 U1518 ( .A(n1593), .B(n1594), .Y(n1408) );
  OR2X4 U1519 ( .A(n1595), .B(n1596), .Y(n1594) );
  AND2X4 U1520 ( .A(n1597), .B(n1598), .Y(n1593) );
  OR2X4 U1521 ( .A(n1402), .B(n1404), .Y(n1406) );
  AND2X4 U1522 ( .A(n1599), .B(n1217), .Y(Y[17]) );
  OR2X4 U1523 ( .A(n1600), .B(n1601), .Y(n1217) );
  OR2X4 U1524 ( .A(n1602), .B(n1603), .Y(n1601) );
  OR2X4 U1525 ( .A(n1604), .B(n1605), .Y(n1599) );
  INVX4 U1526 ( .A(n1603), .Y(n1605) );
  OR2X4 U1527 ( .A(n1606), .B(n1607), .Y(n1603) );
  NOR2X4 U1528 ( .A(n1402), .B(n1404), .Y(n1607) );
  AND2X4 U1529 ( .A(n1404), .B(n1402), .Y(n1606) );
  OR2X4 U1530 ( .A(n1608), .B(n1609), .Y(n1402) );
  OR2X4 U1531 ( .A(n1610), .B(n1611), .Y(n1609) );
  AND2X4 U1532 ( .A(n1612), .B(n1613), .Y(n1611) );
  OR2X4 U1533 ( .A(n1614), .B(n1595), .Y(n1613) );
  NOR2X4 U1534 ( .A(n1615), .B(n1616), .Y(n1595) );
  AND2X4 U1535 ( .A(n1615), .B(n1616), .Y(n1614) );
  AND2X4 U1536 ( .A(n1617), .B(n1597), .Y(n1610) );
  AND2X4 U1537 ( .A(n1616), .B(n1598), .Y(n1617) );
  AND2X4 U1538 ( .A(n1596), .B(n1615), .Y(n1608) );
  INVX4 U1539 ( .A(n1598), .Y(n1615) );
  OR2X4 U1540 ( .A(n1618), .B(n1619), .Y(n1598) );
  AND2X4 U1541 ( .A(n1620), .B(n1621), .Y(n1618) );
  NOR2X4 U1542 ( .A(n1612), .B(n1616), .Y(n1596) );
  OR2X4 U1543 ( .A(n1622), .B(n175), .Y(n1616) );
  INVX4 U1544 ( .A(n1597), .Y(n1612) );
  OR2X4 U1545 ( .A(n1623), .B(n1624), .Y(n1597) );
  AND2X4 U1546 ( .A(n1625), .B(n1626), .Y(n1624) );
  AND2X4 U1547 ( .A(n1627), .B(n1424), .Y(n1626) );
  OR2X4 U1548 ( .A(n1628), .B(n1629), .Y(n1424) );
  OR2X4 U1549 ( .A(n1630), .B(n1631), .Y(n1627) );
  INVX4 U1550 ( .A(n1423), .Y(n1625) );
  AND2X4 U1551 ( .A(n1423), .B(n1632), .Y(n1623) );
  OR2X4 U1552 ( .A(n1633), .B(n1422), .Y(n1632) );
  AND2X4 U1553 ( .A(n1629), .B(n1628), .Y(n1422) );
  AND2X4 U1554 ( .A(n1630), .B(n1631), .Y(n1633) );
  INVX4 U1555 ( .A(n1628), .Y(n1631) );
  AND2X4 U1556 ( .A(B[3]), .B(A[14]), .Y(n1628) );
  INVX4 U1557 ( .A(n1629), .Y(n1630) );
  OR2X4 U1558 ( .A(n1634), .B(n1635), .Y(n1629) );
  AND2X4 U1559 ( .A(n1636), .B(n1637), .Y(n1634) );
  OR2X4 U1560 ( .A(n1638), .B(n1639), .Y(n1423) );
  AND2X4 U1561 ( .A(n1640), .B(n1641), .Y(n1639) );
  AND2X4 U1562 ( .A(n1642), .B(n1439), .Y(n1641) );
  OR2X4 U1563 ( .A(n1643), .B(n1644), .Y(n1439) );
  OR2X4 U1564 ( .A(n1645), .B(n1646), .Y(n1642) );
  INVX4 U1565 ( .A(n1438), .Y(n1640) );
  AND2X4 U1566 ( .A(n1438), .B(n1647), .Y(n1638) );
  OR2X4 U1567 ( .A(n1648), .B(n1437), .Y(n1647) );
  AND2X4 U1568 ( .A(n1644), .B(n1643), .Y(n1437) );
  AND2X4 U1569 ( .A(n1645), .B(n1646), .Y(n1648) );
  INVX4 U1570 ( .A(n1643), .Y(n1646) );
  AND2X4 U1571 ( .A(B[4]), .B(A[13]), .Y(n1643) );
  INVX4 U1572 ( .A(n1644), .Y(n1645) );
  OR2X4 U1573 ( .A(n1649), .B(n1650), .Y(n1644) );
  AND2X4 U1574 ( .A(n1651), .B(n1652), .Y(n1649) );
  OR2X4 U1575 ( .A(n1653), .B(n1654), .Y(n1438) );
  AND2X4 U1576 ( .A(n1655), .B(n1656), .Y(n1654) );
  AND2X4 U1577 ( .A(n1657), .B(n1454), .Y(n1656) );
  OR2X4 U1578 ( .A(n1658), .B(n1659), .Y(n1454) );
  OR2X4 U1579 ( .A(n1660), .B(n1661), .Y(n1657) );
  INVX4 U1580 ( .A(n1453), .Y(n1655) );
  AND2X4 U1581 ( .A(n1453), .B(n1662), .Y(n1653) );
  OR2X4 U1582 ( .A(n1663), .B(n1452), .Y(n1662) );
  AND2X4 U1583 ( .A(n1659), .B(n1658), .Y(n1452) );
  AND2X4 U1584 ( .A(n1660), .B(n1661), .Y(n1663) );
  INVX4 U1585 ( .A(n1658), .Y(n1661) );
  AND2X4 U1586 ( .A(B[5]), .B(A[12]), .Y(n1658) );
  INVX4 U1587 ( .A(n1659), .Y(n1660) );
  OR2X4 U1588 ( .A(n1664), .B(n1665), .Y(n1659) );
  AND2X4 U1589 ( .A(n1666), .B(n1667), .Y(n1664) );
  OR2X4 U1590 ( .A(n1668), .B(n1669), .Y(n1453) );
  AND2X4 U1591 ( .A(n1670), .B(n1671), .Y(n1669) );
  AND2X4 U1592 ( .A(n1672), .B(n1469), .Y(n1671) );
  OR2X4 U1593 ( .A(n1673), .B(n1674), .Y(n1469) );
  OR2X4 U1594 ( .A(n1675), .B(n1676), .Y(n1672) );
  INVX4 U1595 ( .A(n1468), .Y(n1670) );
  AND2X4 U1596 ( .A(n1468), .B(n1677), .Y(n1668) );
  OR2X4 U1597 ( .A(n1678), .B(n1467), .Y(n1677) );
  AND2X4 U1598 ( .A(n1674), .B(n1673), .Y(n1467) );
  AND2X4 U1599 ( .A(n1675), .B(n1676), .Y(n1678) );
  INVX4 U1600 ( .A(n1673), .Y(n1676) );
  AND2X4 U1601 ( .A(B[6]), .B(A[11]), .Y(n1673) );
  INVX4 U1602 ( .A(n1674), .Y(n1675) );
  OR2X4 U1603 ( .A(n1679), .B(n1680), .Y(n1674) );
  AND2X4 U1604 ( .A(n1681), .B(n1682), .Y(n1679) );
  OR2X4 U1605 ( .A(n1683), .B(n1684), .Y(n1468) );
  AND2X4 U1606 ( .A(n1685), .B(n1686), .Y(n1684) );
  AND2X4 U1607 ( .A(n1687), .B(n1484), .Y(n1686) );
  OR2X4 U1608 ( .A(n1688), .B(n1689), .Y(n1484) );
  OR2X4 U1609 ( .A(n1690), .B(n1691), .Y(n1687) );
  INVX4 U1610 ( .A(n1483), .Y(n1685) );
  AND2X4 U1611 ( .A(n1483), .B(n1692), .Y(n1683) );
  OR2X4 U1612 ( .A(n1693), .B(n1482), .Y(n1692) );
  AND2X4 U1613 ( .A(n1689), .B(n1688), .Y(n1482) );
  AND2X4 U1614 ( .A(n1690), .B(n1691), .Y(n1693) );
  INVX4 U1615 ( .A(n1688), .Y(n1691) );
  AND2X4 U1616 ( .A(B[7]), .B(A[10]), .Y(n1688) );
  INVX4 U1617 ( .A(n1689), .Y(n1690) );
  OR2X4 U1618 ( .A(n1694), .B(n1695), .Y(n1689) );
  AND2X4 U1619 ( .A(n1696), .B(n1697), .Y(n1694) );
  OR2X4 U1620 ( .A(n1698), .B(n1699), .Y(n1483) );
  AND2X4 U1621 ( .A(n1700), .B(n1701), .Y(n1699) );
  AND2X4 U1622 ( .A(n1702), .B(n1499), .Y(n1701) );
  OR2X4 U1623 ( .A(n1703), .B(n1704), .Y(n1499) );
  OR2X4 U1624 ( .A(n1705), .B(n1706), .Y(n1702) );
  INVX4 U1625 ( .A(n1498), .Y(n1700) );
  AND2X4 U1626 ( .A(n1498), .B(n1707), .Y(n1698) );
  OR2X4 U1627 ( .A(n1708), .B(n1497), .Y(n1707) );
  AND2X4 U1628 ( .A(n1704), .B(n1703), .Y(n1497) );
  AND2X4 U1629 ( .A(n1705), .B(n1706), .Y(n1708) );
  INVX4 U1630 ( .A(n1703), .Y(n1706) );
  AND2X4 U1631 ( .A(B[8]), .B(A[9]), .Y(n1703) );
  INVX4 U1632 ( .A(n1704), .Y(n1705) );
  OR2X4 U1633 ( .A(n1709), .B(n1710), .Y(n1704) );
  AND2X4 U1634 ( .A(n1711), .B(n1712), .Y(n1709) );
  OR2X4 U1635 ( .A(n1713), .B(n1714), .Y(n1498) );
  AND2X4 U1636 ( .A(n1715), .B(n1716), .Y(n1714) );
  AND2X4 U1637 ( .A(n1717), .B(n1514), .Y(n1716) );
  OR2X4 U1638 ( .A(n1718), .B(n1719), .Y(n1514) );
  OR2X4 U1639 ( .A(n1720), .B(n1721), .Y(n1717) );
  INVX4 U1640 ( .A(n1513), .Y(n1715) );
  AND2X4 U1641 ( .A(n1513), .B(n1722), .Y(n1713) );
  OR2X4 U1642 ( .A(n1723), .B(n1512), .Y(n1722) );
  AND2X4 U1643 ( .A(n1719), .B(n1718), .Y(n1512) );
  AND2X4 U1644 ( .A(n1720), .B(n1721), .Y(n1723) );
  INVX4 U1645 ( .A(n1718), .Y(n1721) );
  AND2X4 U1646 ( .A(B[9]), .B(A[8]), .Y(n1718) );
  INVX4 U1647 ( .A(n1719), .Y(n1720) );
  OR2X4 U1648 ( .A(n1724), .B(n1725), .Y(n1719) );
  AND2X4 U1649 ( .A(n1726), .B(n1727), .Y(n1724) );
  OR2X4 U1650 ( .A(n1728), .B(n1729), .Y(n1513) );
  AND2X4 U1651 ( .A(n1730), .B(n1731), .Y(n1729) );
  AND2X4 U1652 ( .A(n1732), .B(n1529), .Y(n1731) );
  OR2X4 U1653 ( .A(n1733), .B(n1734), .Y(n1529) );
  OR2X4 U1654 ( .A(n1735), .B(n1736), .Y(n1732) );
  INVX4 U1655 ( .A(n1528), .Y(n1730) );
  AND2X4 U1656 ( .A(n1528), .B(n1737), .Y(n1728) );
  OR2X4 U1657 ( .A(n1738), .B(n1527), .Y(n1737) );
  AND2X4 U1658 ( .A(n1734), .B(n1733), .Y(n1527) );
  AND2X4 U1659 ( .A(n1735), .B(n1736), .Y(n1738) );
  INVX4 U1660 ( .A(n1733), .Y(n1736) );
  AND2X4 U1661 ( .A(A[7]), .B(B[10]), .Y(n1733) );
  INVX4 U1662 ( .A(n1734), .Y(n1735) );
  OR2X4 U1663 ( .A(n1739), .B(n1740), .Y(n1734) );
  AND2X4 U1664 ( .A(n1741), .B(n1742), .Y(n1739) );
  OR2X4 U1665 ( .A(n1743), .B(n1744), .Y(n1528) );
  AND2X4 U1666 ( .A(n1745), .B(n1746), .Y(n1744) );
  AND2X4 U1667 ( .A(n1747), .B(n1544), .Y(n1746) );
  OR2X4 U1668 ( .A(n1748), .B(n1749), .Y(n1544) );
  OR2X4 U1669 ( .A(n1750), .B(n1751), .Y(n1747) );
  INVX4 U1670 ( .A(n1543), .Y(n1745) );
  AND2X4 U1671 ( .A(n1543), .B(n1752), .Y(n1743) );
  OR2X4 U1672 ( .A(n1753), .B(n1542), .Y(n1752) );
  AND2X4 U1673 ( .A(n1749), .B(n1748), .Y(n1542) );
  AND2X4 U1674 ( .A(n1750), .B(n1751), .Y(n1753) );
  INVX4 U1675 ( .A(n1748), .Y(n1751) );
  AND2X4 U1676 ( .A(A[6]), .B(B[11]), .Y(n1748) );
  INVX4 U1677 ( .A(n1749), .Y(n1750) );
  OR2X4 U1678 ( .A(n1754), .B(n1755), .Y(n1749) );
  AND2X4 U1679 ( .A(n1756), .B(n1757), .Y(n1754) );
  OR2X4 U1680 ( .A(n1758), .B(n1759), .Y(n1543) );
  AND2X4 U1681 ( .A(n1760), .B(n1761), .Y(n1759) );
  AND2X4 U1682 ( .A(n1762), .B(n1559), .Y(n1761) );
  OR2X4 U1683 ( .A(n1763), .B(n1764), .Y(n1559) );
  OR2X4 U1684 ( .A(n1765), .B(n1766), .Y(n1762) );
  INVX4 U1685 ( .A(n1558), .Y(n1760) );
  AND2X4 U1686 ( .A(n1558), .B(n1767), .Y(n1758) );
  OR2X4 U1687 ( .A(n1768), .B(n1557), .Y(n1767) );
  AND2X4 U1688 ( .A(n1764), .B(n1763), .Y(n1557) );
  AND2X4 U1689 ( .A(n1765), .B(n1766), .Y(n1768) );
  INVX4 U1690 ( .A(n1763), .Y(n1766) );
  AND2X4 U1691 ( .A(A[5]), .B(B[12]), .Y(n1763) );
  INVX4 U1692 ( .A(n1764), .Y(n1765) );
  OR2X4 U1693 ( .A(n1769), .B(n1770), .Y(n1764) );
  AND2X4 U1694 ( .A(n1771), .B(n1772), .Y(n1769) );
  OR2X4 U1695 ( .A(n1773), .B(n1774), .Y(n1558) );
  AND2X4 U1696 ( .A(n1775), .B(n1776), .Y(n1774) );
  AND2X4 U1697 ( .A(n1777), .B(n1574), .Y(n1776) );
  OR2X4 U1698 ( .A(n1778), .B(n1779), .Y(n1574) );
  OR2X4 U1699 ( .A(n1780), .B(n1781), .Y(n1777) );
  INVX4 U1700 ( .A(n1573), .Y(n1775) );
  AND2X4 U1701 ( .A(n1573), .B(n1782), .Y(n1773) );
  OR2X4 U1702 ( .A(n1783), .B(n1572), .Y(n1782) );
  AND2X4 U1703 ( .A(n1779), .B(n1778), .Y(n1572) );
  AND2X4 U1704 ( .A(n1780), .B(n1781), .Y(n1783) );
  INVX4 U1705 ( .A(n1778), .Y(n1781) );
  AND2X4 U1706 ( .A(A[4]), .B(B[13]), .Y(n1778) );
  INVX4 U1707 ( .A(n1779), .Y(n1780) );
  OR2X4 U1708 ( .A(n1784), .B(n1785), .Y(n1779) );
  AND2X4 U1709 ( .A(n1786), .B(n1787), .Y(n1784) );
  OR2X4 U1710 ( .A(n1788), .B(n1789), .Y(n1786) );
  OR2X4 U1711 ( .A(n1790), .B(n1791), .Y(n1573) );
  AND2X4 U1712 ( .A(n1792), .B(n1793), .Y(n1791) );
  INVX4 U1713 ( .A(n1589), .Y(n1793) );
  OR2X4 U1714 ( .A(n1794), .B(n1795), .Y(n1792) );
  AND2X4 U1715 ( .A(A[3]), .B(n1796), .Y(n1795) );
  OR2X4 U1716 ( .A(n1797), .B(n293), .Y(n1796) );
  AND2X4 U1717 ( .A(B[14]), .B(n142), .Y(n1797) );
  AND2X4 U1718 ( .A(A[2]), .B(n1798), .Y(n1794) );
  OR2X4 U1719 ( .A(n1799), .B(n297), .Y(n1798) );
  AND2X4 U1720 ( .A(B[15]), .B(n1583), .Y(n1799) );
  AND2X4 U1721 ( .A(n1589), .B(n1800), .Y(n1790) );
  OR2X4 U1722 ( .A(n1588), .B(n1801), .Y(n1800) );
  AND2X4 U1723 ( .A(n142), .B(n1583), .Y(n1801) );
  INVX4 U1724 ( .A(A[3]), .Y(n1583) );
  AND2X4 U1725 ( .A(n1802), .B(n306), .Y(n1588) );
  AND2X4 U1726 ( .A(A[3]), .B(A[2]), .Y(n1802) );
  AND2X4 U1727 ( .A(n1803), .B(n306), .Y(n1589) );
  AND2X4 U1728 ( .A(B[14]), .B(B[15]), .Y(n306) );
  NAND2X4 U1729 ( .A(n1804), .B(n1805), .Y(n1803) );
  OR2X4 U1730 ( .A(n1806), .B(n142), .Y(n1805) );
  NOR2X4 U1731 ( .A(n1807), .B(n1808), .Y(n1404) );
  OR2X4 U1732 ( .A(n1809), .B(n1810), .Y(n1808) );
  AND2X4 U1733 ( .A(n1811), .B(n1812), .Y(n1807) );
  AND2X4 U1734 ( .A(n1813), .B(n1814), .Y(n1604) );
  AND2X4 U1735 ( .A(n1815), .B(n1816), .Y(Y[16]) );
  OR2X4 U1736 ( .A(n1602), .B(n1600), .Y(n1816) );
  INVX4 U1737 ( .A(n1814), .Y(n1602) );
  OR2X4 U1738 ( .A(n1813), .B(n1814), .Y(n1815) );
  OR2X4 U1739 ( .A(n1817), .B(n1818), .Y(n1814) );
  AND2X4 U1740 ( .A(n1819), .B(n1820), .Y(n1817) );
  INVX4 U1741 ( .A(n1600), .Y(n1813) );
  OR2X4 U1742 ( .A(n1821), .B(n1822), .Y(n1600) );
  OR2X4 U1743 ( .A(n1823), .B(n1824), .Y(n1822) );
  AND2X4 U1744 ( .A(n1825), .B(n1826), .Y(n1824) );
  OR2X4 U1745 ( .A(n1827), .B(n1809), .Y(n1826) );
  NOR2X4 U1746 ( .A(n1828), .B(n1829), .Y(n1809) );
  AND2X4 U1747 ( .A(n1828), .B(n1829), .Y(n1827) );
  AND2X4 U1748 ( .A(n1830), .B(n1811), .Y(n1823) );
  AND2X4 U1749 ( .A(n1829), .B(n1812), .Y(n1830) );
  AND2X4 U1750 ( .A(n1810), .B(n1828), .Y(n1821) );
  INVX4 U1751 ( .A(n1812), .Y(n1828) );
  OR2X4 U1752 ( .A(n1831), .B(n1832), .Y(n1812) );
  AND2X4 U1753 ( .A(n1833), .B(n1834), .Y(n1831) );
  NOR2X4 U1754 ( .A(n1825), .B(n1829), .Y(n1810) );
  OR2X4 U1755 ( .A(n132), .B(n175), .Y(n1829) );
  INVX4 U1756 ( .A(A[15]), .Y(n175) );
  INVX4 U1757 ( .A(n1811), .Y(n1825) );
  OR2X4 U1758 ( .A(n1835), .B(n1836), .Y(n1811) );
  AND2X4 U1759 ( .A(n1837), .B(n1838), .Y(n1836) );
  AND2X4 U1760 ( .A(n1839), .B(n1621), .Y(n1838) );
  OR2X4 U1761 ( .A(n1840), .B(n1841), .Y(n1621) );
  OR2X4 U1762 ( .A(n1842), .B(n1843), .Y(n1839) );
  INVX4 U1763 ( .A(n1620), .Y(n1837) );
  AND2X4 U1764 ( .A(n1620), .B(n1844), .Y(n1835) );
  OR2X4 U1765 ( .A(n1845), .B(n1619), .Y(n1844) );
  AND2X4 U1766 ( .A(n1841), .B(n1840), .Y(n1619) );
  AND2X4 U1767 ( .A(n1842), .B(n1843), .Y(n1845) );
  INVX4 U1768 ( .A(n1840), .Y(n1843) );
  AND2X4 U1769 ( .A(B[2]), .B(A[14]), .Y(n1840) );
  INVX4 U1770 ( .A(n1841), .Y(n1842) );
  OR2X4 U1771 ( .A(n1846), .B(n1847), .Y(n1841) );
  AND2X4 U1772 ( .A(n1848), .B(n1849), .Y(n1846) );
  OR2X4 U1773 ( .A(n1850), .B(n1851), .Y(n1620) );
  AND2X4 U1774 ( .A(n1852), .B(n1853), .Y(n1851) );
  AND2X4 U1775 ( .A(n1854), .B(n1637), .Y(n1853) );
  OR2X4 U1776 ( .A(n1855), .B(n1856), .Y(n1637) );
  OR2X4 U1777 ( .A(n1857), .B(n1858), .Y(n1854) );
  INVX4 U1778 ( .A(n1636), .Y(n1852) );
  AND2X4 U1779 ( .A(n1636), .B(n1859), .Y(n1850) );
  OR2X4 U1780 ( .A(n1860), .B(n1635), .Y(n1859) );
  AND2X4 U1781 ( .A(n1856), .B(n1855), .Y(n1635) );
  AND2X4 U1782 ( .A(n1857), .B(n1858), .Y(n1860) );
  INVX4 U1783 ( .A(n1855), .Y(n1858) );
  AND2X4 U1784 ( .A(B[3]), .B(A[13]), .Y(n1855) );
  INVX4 U1785 ( .A(n1856), .Y(n1857) );
  OR2X4 U1786 ( .A(n1861), .B(n1862), .Y(n1856) );
  AND2X4 U1787 ( .A(n1863), .B(n1864), .Y(n1861) );
  OR2X4 U1788 ( .A(n1865), .B(n1866), .Y(n1636) );
  AND2X4 U1789 ( .A(n1867), .B(n1868), .Y(n1866) );
  AND2X4 U1790 ( .A(n1869), .B(n1652), .Y(n1868) );
  OR2X4 U1791 ( .A(n1870), .B(n1871), .Y(n1652) );
  OR2X4 U1792 ( .A(n1872), .B(n1873), .Y(n1869) );
  INVX4 U1793 ( .A(n1651), .Y(n1867) );
  AND2X4 U1794 ( .A(n1651), .B(n1874), .Y(n1865) );
  OR2X4 U1795 ( .A(n1875), .B(n1650), .Y(n1874) );
  AND2X4 U1796 ( .A(n1871), .B(n1870), .Y(n1650) );
  AND2X4 U1797 ( .A(n1872), .B(n1873), .Y(n1875) );
  INVX4 U1798 ( .A(n1870), .Y(n1873) );
  AND2X4 U1799 ( .A(B[4]), .B(A[12]), .Y(n1870) );
  INVX4 U1800 ( .A(n1871), .Y(n1872) );
  OR2X4 U1801 ( .A(n1876), .B(n1877), .Y(n1871) );
  AND2X4 U1802 ( .A(n1878), .B(n1879), .Y(n1876) );
  OR2X4 U1803 ( .A(n1880), .B(n1881), .Y(n1651) );
  AND2X4 U1804 ( .A(n1882), .B(n1883), .Y(n1881) );
  AND2X4 U1805 ( .A(n1884), .B(n1667), .Y(n1883) );
  OR2X4 U1806 ( .A(n1885), .B(n1886), .Y(n1667) );
  OR2X4 U1807 ( .A(n1887), .B(n1888), .Y(n1884) );
  INVX4 U1808 ( .A(n1666), .Y(n1882) );
  AND2X4 U1809 ( .A(n1666), .B(n1889), .Y(n1880) );
  OR2X4 U1810 ( .A(n1890), .B(n1665), .Y(n1889) );
  AND2X4 U1811 ( .A(n1886), .B(n1885), .Y(n1665) );
  AND2X4 U1812 ( .A(n1887), .B(n1888), .Y(n1890) );
  INVX4 U1813 ( .A(n1885), .Y(n1888) );
  AND2X4 U1814 ( .A(B[5]), .B(A[11]), .Y(n1885) );
  INVX4 U1815 ( .A(n1886), .Y(n1887) );
  OR2X4 U1816 ( .A(n1891), .B(n1892), .Y(n1886) );
  AND2X4 U1817 ( .A(n1893), .B(n1894), .Y(n1891) );
  OR2X4 U1818 ( .A(n1895), .B(n1896), .Y(n1666) );
  AND2X4 U1819 ( .A(n1897), .B(n1898), .Y(n1896) );
  AND2X4 U1820 ( .A(n1899), .B(n1682), .Y(n1898) );
  OR2X4 U1821 ( .A(n1900), .B(n1901), .Y(n1682) );
  OR2X4 U1822 ( .A(n1902), .B(n1903), .Y(n1899) );
  INVX4 U1823 ( .A(n1681), .Y(n1897) );
  AND2X4 U1824 ( .A(n1681), .B(n1904), .Y(n1895) );
  OR2X4 U1825 ( .A(n1905), .B(n1680), .Y(n1904) );
  AND2X4 U1826 ( .A(n1901), .B(n1900), .Y(n1680) );
  AND2X4 U1827 ( .A(n1902), .B(n1903), .Y(n1905) );
  INVX4 U1828 ( .A(n1900), .Y(n1903) );
  AND2X4 U1829 ( .A(B[6]), .B(A[10]), .Y(n1900) );
  INVX4 U1830 ( .A(n1901), .Y(n1902) );
  OR2X4 U1831 ( .A(n1906), .B(n1907), .Y(n1901) );
  AND2X4 U1832 ( .A(n1908), .B(n1909), .Y(n1906) );
  OR2X4 U1833 ( .A(n1910), .B(n1911), .Y(n1681) );
  AND2X4 U1834 ( .A(n1912), .B(n1913), .Y(n1911) );
  AND2X4 U1835 ( .A(n1914), .B(n1697), .Y(n1913) );
  OR2X4 U1836 ( .A(n1915), .B(n1916), .Y(n1697) );
  OR2X4 U1837 ( .A(n1917), .B(n1918), .Y(n1914) );
  INVX4 U1838 ( .A(n1696), .Y(n1912) );
  AND2X4 U1839 ( .A(n1696), .B(n1919), .Y(n1910) );
  OR2X4 U1840 ( .A(n1920), .B(n1695), .Y(n1919) );
  AND2X4 U1841 ( .A(n1916), .B(n1915), .Y(n1695) );
  AND2X4 U1842 ( .A(n1917), .B(n1918), .Y(n1920) );
  INVX4 U1843 ( .A(n1915), .Y(n1918) );
  AND2X4 U1844 ( .A(B[7]), .B(A[9]), .Y(n1915) );
  INVX4 U1845 ( .A(n1916), .Y(n1917) );
  OR2X4 U1846 ( .A(n1921), .B(n1922), .Y(n1916) );
  AND2X4 U1847 ( .A(n1923), .B(n1924), .Y(n1921) );
  OR2X4 U1848 ( .A(n1925), .B(n1926), .Y(n1696) );
  AND2X4 U1849 ( .A(n1927), .B(n1928), .Y(n1926) );
  AND2X4 U1850 ( .A(n1929), .B(n1712), .Y(n1928) );
  OR2X4 U1851 ( .A(n1930), .B(n1931), .Y(n1712) );
  OR2X4 U1852 ( .A(n1932), .B(n1933), .Y(n1929) );
  INVX4 U1853 ( .A(n1711), .Y(n1927) );
  AND2X4 U1854 ( .A(n1711), .B(n1934), .Y(n1925) );
  OR2X4 U1855 ( .A(n1935), .B(n1710), .Y(n1934) );
  AND2X4 U1856 ( .A(n1931), .B(n1930), .Y(n1710) );
  AND2X4 U1857 ( .A(n1932), .B(n1933), .Y(n1935) );
  INVX4 U1858 ( .A(n1930), .Y(n1933) );
  AND2X4 U1859 ( .A(B[8]), .B(A[8]), .Y(n1930) );
  INVX4 U1860 ( .A(n1931), .Y(n1932) );
  OR2X4 U1861 ( .A(n1936), .B(n1937), .Y(n1931) );
  AND2X4 U1862 ( .A(n1938), .B(n1939), .Y(n1936) );
  OR2X4 U1863 ( .A(n1940), .B(n1941), .Y(n1711) );
  AND2X4 U1864 ( .A(n1942), .B(n1943), .Y(n1941) );
  AND2X4 U1865 ( .A(n1944), .B(n1727), .Y(n1943) );
  OR2X4 U1866 ( .A(n1945), .B(n1946), .Y(n1727) );
  OR2X4 U1867 ( .A(n1947), .B(n1948), .Y(n1944) );
  INVX4 U1868 ( .A(n1726), .Y(n1942) );
  AND2X4 U1869 ( .A(n1726), .B(n1949), .Y(n1940) );
  OR2X4 U1870 ( .A(n1950), .B(n1725), .Y(n1949) );
  AND2X4 U1871 ( .A(n1946), .B(n1945), .Y(n1725) );
  AND2X4 U1872 ( .A(n1947), .B(n1948), .Y(n1950) );
  INVX4 U1873 ( .A(n1945), .Y(n1948) );
  AND2X4 U1874 ( .A(B[9]), .B(A[7]), .Y(n1945) );
  INVX4 U1875 ( .A(n1946), .Y(n1947) );
  OR2X4 U1876 ( .A(n1951), .B(n1952), .Y(n1946) );
  AND2X4 U1877 ( .A(n1953), .B(n1954), .Y(n1951) );
  OR2X4 U1878 ( .A(n1955), .B(n1956), .Y(n1726) );
  AND2X4 U1879 ( .A(n1957), .B(n1958), .Y(n1956) );
  AND2X4 U1880 ( .A(n1959), .B(n1742), .Y(n1958) );
  OR2X4 U1881 ( .A(n1960), .B(n1961), .Y(n1742) );
  OR2X4 U1882 ( .A(n1962), .B(n1963), .Y(n1959) );
  INVX4 U1883 ( .A(n1741), .Y(n1957) );
  AND2X4 U1884 ( .A(n1741), .B(n1964), .Y(n1955) );
  OR2X4 U1885 ( .A(n1965), .B(n1740), .Y(n1964) );
  AND2X4 U1886 ( .A(n1961), .B(n1960), .Y(n1740) );
  AND2X4 U1887 ( .A(n1962), .B(n1963), .Y(n1965) );
  INVX4 U1888 ( .A(n1960), .Y(n1963) );
  AND2X4 U1889 ( .A(A[6]), .B(B[10]), .Y(n1960) );
  INVX4 U1890 ( .A(n1961), .Y(n1962) );
  OR2X4 U1891 ( .A(n1966), .B(n1967), .Y(n1961) );
  AND2X4 U1892 ( .A(n1968), .B(n1969), .Y(n1966) );
  OR2X4 U1893 ( .A(n1970), .B(n1971), .Y(n1741) );
  AND2X4 U1894 ( .A(n1972), .B(n1973), .Y(n1971) );
  AND2X4 U1895 ( .A(n1974), .B(n1757), .Y(n1973) );
  OR2X4 U1896 ( .A(n1975), .B(n1976), .Y(n1757) );
  OR2X4 U1897 ( .A(n1977), .B(n1978), .Y(n1974) );
  INVX4 U1898 ( .A(n1756), .Y(n1972) );
  AND2X4 U1899 ( .A(n1756), .B(n1979), .Y(n1970) );
  OR2X4 U1900 ( .A(n1980), .B(n1755), .Y(n1979) );
  AND2X4 U1901 ( .A(n1976), .B(n1975), .Y(n1755) );
  AND2X4 U1902 ( .A(n1977), .B(n1978), .Y(n1980) );
  INVX4 U1903 ( .A(n1975), .Y(n1978) );
  AND2X4 U1904 ( .A(A[5]), .B(B[11]), .Y(n1975) );
  INVX4 U1905 ( .A(n1976), .Y(n1977) );
  OR2X4 U1906 ( .A(n1981), .B(n1982), .Y(n1976) );
  AND2X4 U1907 ( .A(n1983), .B(n1984), .Y(n1981) );
  OR2X4 U1908 ( .A(n1985), .B(n1986), .Y(n1756) );
  AND2X4 U1909 ( .A(n1987), .B(n1988), .Y(n1986) );
  AND2X4 U1910 ( .A(n1989), .B(n1772), .Y(n1988) );
  OR2X4 U1911 ( .A(n1990), .B(n1991), .Y(n1772) );
  OR2X4 U1912 ( .A(n1992), .B(n1993), .Y(n1989) );
  INVX4 U1913 ( .A(n1771), .Y(n1987) );
  AND2X4 U1914 ( .A(n1771), .B(n1994), .Y(n1985) );
  OR2X4 U1915 ( .A(n1995), .B(n1770), .Y(n1994) );
  AND2X4 U1916 ( .A(n1991), .B(n1990), .Y(n1770) );
  AND2X4 U1917 ( .A(n1992), .B(n1993), .Y(n1995) );
  INVX4 U1918 ( .A(n1990), .Y(n1993) );
  AND2X4 U1919 ( .A(A[4]), .B(B[12]), .Y(n1990) );
  INVX4 U1920 ( .A(n1991), .Y(n1992) );
  OR2X4 U1921 ( .A(n1996), .B(n1997), .Y(n1991) );
  AND2X4 U1922 ( .A(n1998), .B(n1999), .Y(n1996) );
  OR2X4 U1923 ( .A(n2000), .B(n2001), .Y(n1999) );
  OR2X4 U1924 ( .A(n2002), .B(n2003), .Y(n1771) );
  AND2X4 U1925 ( .A(n2004), .B(n2005), .Y(n2003) );
  OR2X4 U1926 ( .A(n2006), .B(n2007), .Y(n2005) );
  AND2X4 U1927 ( .A(n1788), .B(n2008), .Y(n2007) );
  AND2X4 U1928 ( .A(n1789), .B(n2009), .Y(n2006) );
  INVX4 U1929 ( .A(n1787), .Y(n2004) );
  AND2X4 U1930 ( .A(n2010), .B(n1787), .Y(n2002) );
  OR2X4 U1931 ( .A(n2011), .B(n2012), .Y(n1787) );
  OR2X4 U1932 ( .A(n2013), .B(n2014), .Y(n2012) );
  AND2X4 U1933 ( .A(n2015), .B(n142), .Y(n2014) );
  AND2X4 U1934 ( .A(B[15]), .B(n1210), .Y(n2015) );
  AND2X4 U1935 ( .A(A[2]), .B(n2016), .Y(n2013) );
  OR2X4 U1936 ( .A(n2017), .B(n293), .Y(n2016) );
  NOR2X4 U1937 ( .A(n183), .B(n1210), .Y(n2017) );
  AND2X4 U1938 ( .A(n297), .B(A[1]), .Y(n2011) );
  OR2X4 U1939 ( .A(n2018), .B(n1785), .Y(n2010) );
  AND2X4 U1940 ( .A(n1789), .B(n1788), .Y(n1785) );
  INVX4 U1941 ( .A(n2008), .Y(n1789) );
  AND2X4 U1942 ( .A(n2009), .B(n2008), .Y(n2018) );
  OR2X4 U1943 ( .A(n2019), .B(n2020), .Y(n2008) );
  AND2X4 U1944 ( .A(n2021), .B(n2022), .Y(n2019) );
  OR2X4 U1945 ( .A(n2023), .B(n183), .Y(n2022) );
  AND2X4 U1946 ( .A(n2024), .B(n2025), .Y(n2023) );
  OR2X4 U1947 ( .A(n2026), .B(n1804), .Y(n2025) );
  OR2X4 U1948 ( .A(n2026), .B(n142), .Y(n2021) );
  INVX4 U1949 ( .A(n1788), .Y(n2009) );
  AND2X4 U1950 ( .A(A[3]), .B(B[13]), .Y(n1788) );
  OR2X4 U1951 ( .A(n2027), .B(n2028), .Y(Y[15]) );
  AND2X4 U1952 ( .A(n2029), .B(n2030), .Y(n2028) );
  AND2X4 U1953 ( .A(n2031), .B(n1820), .Y(n2030) );
  OR2X4 U1954 ( .A(n2032), .B(n2033), .Y(n1820) );
  OR2X4 U1955 ( .A(n2034), .B(n2035), .Y(n2031) );
  INVX4 U1956 ( .A(n1819), .Y(n2029) );
  AND2X4 U1957 ( .A(n1819), .B(n2036), .Y(n2027) );
  OR2X4 U1958 ( .A(n2037), .B(n1818), .Y(n2036) );
  AND2X4 U1959 ( .A(n2033), .B(n2032), .Y(n1818) );
  AND2X4 U1960 ( .A(n2034), .B(n2035), .Y(n2037) );
  INVX4 U1961 ( .A(n2032), .Y(n2035) );
  AND2X4 U1962 ( .A(B[0]), .B(A[15]), .Y(n2032) );
  INVX4 U1963 ( .A(n2033), .Y(n2034) );
  OR2X4 U1964 ( .A(n2038), .B(n2039), .Y(n2033) );
  AND2X4 U1965 ( .A(n2040), .B(n2041), .Y(n2038) );
  OR2X4 U1966 ( .A(n2042), .B(n2043), .Y(n1819) );
  AND2X4 U1967 ( .A(n2044), .B(n2045), .Y(n2043) );
  AND2X4 U1968 ( .A(n2046), .B(n1834), .Y(n2045) );
  OR2X4 U1969 ( .A(n2047), .B(n2048), .Y(n1834) );
  OR2X4 U1970 ( .A(n2049), .B(n2050), .Y(n2046) );
  INVX4 U1971 ( .A(n1833), .Y(n2044) );
  AND2X4 U1972 ( .A(n1833), .B(n2051), .Y(n2042) );
  OR2X4 U1973 ( .A(n2052), .B(n1832), .Y(n2051) );
  AND2X4 U1974 ( .A(n2048), .B(n2047), .Y(n1832) );
  AND2X4 U1975 ( .A(n2049), .B(n2050), .Y(n2052) );
  INVX4 U1976 ( .A(n2047), .Y(n2050) );
  AND2X4 U1977 ( .A(B[1]), .B(A[14]), .Y(n2047) );
  INVX4 U1978 ( .A(n2048), .Y(n2049) );
  OR2X4 U1979 ( .A(n2053), .B(n2054), .Y(n2048) );
  AND2X4 U1980 ( .A(n2055), .B(n2056), .Y(n2053) );
  OR2X4 U1981 ( .A(n2057), .B(n2058), .Y(n1833) );
  AND2X4 U1982 ( .A(n2059), .B(n2060), .Y(n2058) );
  AND2X4 U1983 ( .A(n2061), .B(n1849), .Y(n2060) );
  OR2X4 U1984 ( .A(n2062), .B(n2063), .Y(n1849) );
  OR2X4 U1985 ( .A(n2064), .B(n2065), .Y(n2061) );
  INVX4 U1986 ( .A(n1848), .Y(n2059) );
  AND2X4 U1987 ( .A(n1848), .B(n2066), .Y(n2057) );
  OR2X4 U1988 ( .A(n2067), .B(n1847), .Y(n2066) );
  AND2X4 U1989 ( .A(n2063), .B(n2062), .Y(n1847) );
  AND2X4 U1990 ( .A(n2064), .B(n2065), .Y(n2067) );
  INVX4 U1991 ( .A(n2062), .Y(n2065) );
  AND2X4 U1992 ( .A(B[2]), .B(A[13]), .Y(n2062) );
  INVX4 U1993 ( .A(n2063), .Y(n2064) );
  OR2X4 U1994 ( .A(n2068), .B(n2069), .Y(n2063) );
  AND2X4 U1995 ( .A(n2070), .B(n2071), .Y(n2068) );
  OR2X4 U1996 ( .A(n2072), .B(n2073), .Y(n1848) );
  AND2X4 U1997 ( .A(n2074), .B(n2075), .Y(n2073) );
  AND2X4 U1998 ( .A(n2076), .B(n1864), .Y(n2075) );
  OR2X4 U1999 ( .A(n2077), .B(n2078), .Y(n1864) );
  OR2X4 U2000 ( .A(n2079), .B(n2080), .Y(n2076) );
  INVX4 U2001 ( .A(n1863), .Y(n2074) );
  AND2X4 U2002 ( .A(n1863), .B(n2081), .Y(n2072) );
  OR2X4 U2003 ( .A(n2082), .B(n1862), .Y(n2081) );
  AND2X4 U2004 ( .A(n2078), .B(n2077), .Y(n1862) );
  AND2X4 U2005 ( .A(n2079), .B(n2080), .Y(n2082) );
  INVX4 U2006 ( .A(n2077), .Y(n2080) );
  AND2X4 U2007 ( .A(B[3]), .B(A[12]), .Y(n2077) );
  INVX4 U2008 ( .A(n2078), .Y(n2079) );
  OR2X4 U2009 ( .A(n2083), .B(n2084), .Y(n2078) );
  AND2X4 U2010 ( .A(n2085), .B(n2086), .Y(n2083) );
  OR2X4 U2011 ( .A(n2087), .B(n2088), .Y(n1863) );
  AND2X4 U2012 ( .A(n2089), .B(n2090), .Y(n2088) );
  AND2X4 U2013 ( .A(n2091), .B(n1879), .Y(n2090) );
  OR2X4 U2014 ( .A(n2092), .B(n2093), .Y(n1879) );
  OR2X4 U2015 ( .A(n2094), .B(n2095), .Y(n2091) );
  INVX4 U2016 ( .A(n1878), .Y(n2089) );
  AND2X4 U2017 ( .A(n1878), .B(n2096), .Y(n2087) );
  OR2X4 U2018 ( .A(n2097), .B(n1877), .Y(n2096) );
  AND2X4 U2019 ( .A(n2093), .B(n2092), .Y(n1877) );
  AND2X4 U2020 ( .A(n2094), .B(n2095), .Y(n2097) );
  INVX4 U2021 ( .A(n2092), .Y(n2095) );
  AND2X4 U2022 ( .A(B[4]), .B(A[11]), .Y(n2092) );
  INVX4 U2023 ( .A(n2093), .Y(n2094) );
  OR2X4 U2024 ( .A(n2098), .B(n2099), .Y(n2093) );
  AND2X4 U2025 ( .A(n2100), .B(n2101), .Y(n2098) );
  OR2X4 U2026 ( .A(n2102), .B(n2103), .Y(n1878) );
  AND2X4 U2027 ( .A(n2104), .B(n2105), .Y(n2103) );
  AND2X4 U2028 ( .A(n2106), .B(n1894), .Y(n2105) );
  OR2X4 U2029 ( .A(n2107), .B(n2108), .Y(n1894) );
  OR2X4 U2030 ( .A(n2109), .B(n2110), .Y(n2106) );
  INVX4 U2031 ( .A(n1893), .Y(n2104) );
  AND2X4 U2032 ( .A(n1893), .B(n2111), .Y(n2102) );
  OR2X4 U2033 ( .A(n2112), .B(n1892), .Y(n2111) );
  AND2X4 U2034 ( .A(n2108), .B(n2107), .Y(n1892) );
  AND2X4 U2035 ( .A(n2109), .B(n2110), .Y(n2112) );
  INVX4 U2036 ( .A(n2107), .Y(n2110) );
  AND2X4 U2037 ( .A(B[5]), .B(A[10]), .Y(n2107) );
  INVX4 U2038 ( .A(n2108), .Y(n2109) );
  OR2X4 U2039 ( .A(n2113), .B(n2114), .Y(n2108) );
  AND2X4 U2040 ( .A(n2115), .B(n2116), .Y(n2113) );
  OR2X4 U2041 ( .A(n2117), .B(n2118), .Y(n1893) );
  AND2X4 U2042 ( .A(n2119), .B(n2120), .Y(n2118) );
  AND2X4 U2043 ( .A(n2121), .B(n1909), .Y(n2120) );
  OR2X4 U2044 ( .A(n2122), .B(n2123), .Y(n1909) );
  OR2X4 U2045 ( .A(n2124), .B(n2125), .Y(n2121) );
  INVX4 U2046 ( .A(n1908), .Y(n2119) );
  AND2X4 U2047 ( .A(n1908), .B(n2126), .Y(n2117) );
  OR2X4 U2048 ( .A(n2127), .B(n1907), .Y(n2126) );
  AND2X4 U2049 ( .A(n2123), .B(n2122), .Y(n1907) );
  AND2X4 U2050 ( .A(n2124), .B(n2125), .Y(n2127) );
  INVX4 U2051 ( .A(n2122), .Y(n2125) );
  AND2X4 U2052 ( .A(B[6]), .B(A[9]), .Y(n2122) );
  INVX4 U2053 ( .A(n2123), .Y(n2124) );
  OR2X4 U2054 ( .A(n2128), .B(n2129), .Y(n2123) );
  AND2X4 U2055 ( .A(n2130), .B(n2131), .Y(n2128) );
  OR2X4 U2056 ( .A(n2132), .B(n2133), .Y(n1908) );
  AND2X4 U2057 ( .A(n2134), .B(n2135), .Y(n2133) );
  AND2X4 U2058 ( .A(n2136), .B(n1924), .Y(n2135) );
  OR2X4 U2059 ( .A(n2137), .B(n2138), .Y(n1924) );
  OR2X4 U2060 ( .A(n2139), .B(n2140), .Y(n2136) );
  INVX4 U2061 ( .A(n1923), .Y(n2134) );
  AND2X4 U2062 ( .A(n1923), .B(n2141), .Y(n2132) );
  OR2X4 U2063 ( .A(n2142), .B(n1922), .Y(n2141) );
  AND2X4 U2064 ( .A(n2138), .B(n2137), .Y(n1922) );
  AND2X4 U2065 ( .A(n2139), .B(n2140), .Y(n2142) );
  INVX4 U2066 ( .A(n2137), .Y(n2140) );
  AND2X4 U2067 ( .A(B[7]), .B(A[8]), .Y(n2137) );
  INVX4 U2068 ( .A(n2138), .Y(n2139) );
  OR2X4 U2069 ( .A(n2143), .B(n2144), .Y(n2138) );
  AND2X4 U2070 ( .A(n2145), .B(n2146), .Y(n2143) );
  OR2X4 U2071 ( .A(n2147), .B(n2148), .Y(n1923) );
  AND2X4 U2072 ( .A(n2149), .B(n2150), .Y(n2148) );
  AND2X4 U2073 ( .A(n2151), .B(n1939), .Y(n2150) );
  OR2X4 U2074 ( .A(n2152), .B(n2153), .Y(n1939) );
  OR2X4 U2075 ( .A(n2154), .B(n2155), .Y(n2151) );
  INVX4 U2076 ( .A(n1938), .Y(n2149) );
  AND2X4 U2077 ( .A(n1938), .B(n2156), .Y(n2147) );
  OR2X4 U2078 ( .A(n2157), .B(n1937), .Y(n2156) );
  AND2X4 U2079 ( .A(n2153), .B(n2152), .Y(n1937) );
  AND2X4 U2080 ( .A(n2154), .B(n2155), .Y(n2157) );
  INVX4 U2081 ( .A(n2152), .Y(n2155) );
  AND2X4 U2082 ( .A(B[8]), .B(A[7]), .Y(n2152) );
  INVX4 U2083 ( .A(n2153), .Y(n2154) );
  OR2X4 U2084 ( .A(n2158), .B(n2159), .Y(n2153) );
  AND2X4 U2085 ( .A(n2160), .B(n2161), .Y(n2158) );
  OR2X4 U2086 ( .A(n2162), .B(n2163), .Y(n1938) );
  AND2X4 U2087 ( .A(n2164), .B(n2165), .Y(n2163) );
  AND2X4 U2088 ( .A(n2166), .B(n1954), .Y(n2165) );
  OR2X4 U2089 ( .A(n2167), .B(n2168), .Y(n1954) );
  OR2X4 U2090 ( .A(n2169), .B(n2170), .Y(n2166) );
  INVX4 U2091 ( .A(n1953), .Y(n2164) );
  AND2X4 U2092 ( .A(n1953), .B(n2171), .Y(n2162) );
  OR2X4 U2093 ( .A(n2172), .B(n1952), .Y(n2171) );
  AND2X4 U2094 ( .A(n2168), .B(n2167), .Y(n1952) );
  AND2X4 U2095 ( .A(n2169), .B(n2170), .Y(n2172) );
  INVX4 U2096 ( .A(n2167), .Y(n2170) );
  AND2X4 U2097 ( .A(B[9]), .B(A[6]), .Y(n2167) );
  INVX4 U2098 ( .A(n2168), .Y(n2169) );
  OR2X4 U2099 ( .A(n2173), .B(n2174), .Y(n2168) );
  AND2X4 U2100 ( .A(n2175), .B(n2176), .Y(n2173) );
  OR2X4 U2101 ( .A(n2177), .B(n2178), .Y(n1953) );
  AND2X4 U2102 ( .A(n2179), .B(n2180), .Y(n2178) );
  AND2X4 U2103 ( .A(n2181), .B(n1969), .Y(n2180) );
  OR2X4 U2104 ( .A(n2182), .B(n2183), .Y(n1969) );
  OR2X4 U2105 ( .A(n2184), .B(n2185), .Y(n2181) );
  INVX4 U2106 ( .A(n1968), .Y(n2179) );
  AND2X4 U2107 ( .A(n1968), .B(n2186), .Y(n2177) );
  OR2X4 U2108 ( .A(n2187), .B(n1967), .Y(n2186) );
  AND2X4 U2109 ( .A(n2183), .B(n2182), .Y(n1967) );
  AND2X4 U2110 ( .A(n2184), .B(n2185), .Y(n2187) );
  INVX4 U2111 ( .A(n2182), .Y(n2185) );
  AND2X4 U2112 ( .A(A[5]), .B(B[10]), .Y(n2182) );
  INVX4 U2113 ( .A(n2183), .Y(n2184) );
  OR2X4 U2114 ( .A(n2188), .B(n2189), .Y(n2183) );
  AND2X4 U2115 ( .A(n2190), .B(n2191), .Y(n2188) );
  OR2X4 U2116 ( .A(n2192), .B(n2193), .Y(n1968) );
  AND2X4 U2117 ( .A(n2194), .B(n2195), .Y(n2193) );
  AND2X4 U2118 ( .A(n2196), .B(n1984), .Y(n2195) );
  OR2X4 U2119 ( .A(n2197), .B(n2198), .Y(n1984) );
  OR2X4 U2120 ( .A(n2199), .B(n2200), .Y(n2196) );
  INVX4 U2121 ( .A(n1983), .Y(n2194) );
  AND2X4 U2122 ( .A(n1983), .B(n2201), .Y(n2192) );
  OR2X4 U2123 ( .A(n2202), .B(n1982), .Y(n2201) );
  AND2X4 U2124 ( .A(n2198), .B(n2197), .Y(n1982) );
  AND2X4 U2125 ( .A(n2199), .B(n2200), .Y(n2202) );
  INVX4 U2126 ( .A(n2197), .Y(n2200) );
  AND2X4 U2127 ( .A(A[4]), .B(B[11]), .Y(n2197) );
  INVX4 U2128 ( .A(n2198), .Y(n2199) );
  OR2X4 U2129 ( .A(n2203), .B(n2204), .Y(n2198) );
  AND2X4 U2130 ( .A(n2205), .B(n2206), .Y(n2203) );
  OR2X4 U2131 ( .A(n2207), .B(n2208), .Y(n2206) );
  OR2X4 U2132 ( .A(n2209), .B(n2210), .Y(n1983) );
  AND2X4 U2133 ( .A(n2211), .B(n2212), .Y(n2210) );
  INVX4 U2134 ( .A(n1998), .Y(n2212) );
  OR2X4 U2135 ( .A(n2213), .B(n2214), .Y(n2211) );
  AND2X4 U2136 ( .A(n2000), .B(n2215), .Y(n2214) );
  AND2X4 U2137 ( .A(n2001), .B(n2216), .Y(n2213) );
  AND2X4 U2138 ( .A(n1998), .B(n2217), .Y(n2209) );
  OR2X4 U2139 ( .A(n2218), .B(n1997), .Y(n2217) );
  AND2X4 U2140 ( .A(n2000), .B(n2001), .Y(n1997) );
  INVX4 U2141 ( .A(n2215), .Y(n2001) );
  AND2X4 U2142 ( .A(n2216), .B(n2215), .Y(n2218) );
  OR2X4 U2143 ( .A(n2219), .B(n269), .Y(n2215) );
  AND2X4 U2144 ( .A(n2220), .B(n2221), .Y(n2219) );
  OR2X4 U2145 ( .A(n2222), .B(n2020), .Y(n2221) );
  AND2X4 U2146 ( .A(n2024), .B(n2223), .Y(n2222) );
  OR2X4 U2147 ( .A(n2224), .B(n1804), .Y(n2223) );
  OR2X4 U2148 ( .A(n2224), .B(n142), .Y(n2220) );
  INVX4 U2149 ( .A(n2000), .Y(n2216) );
  AND2X4 U2150 ( .A(A[3]), .B(B[12]), .Y(n2000) );
  OR2X4 U2151 ( .A(n2225), .B(n2226), .Y(n1998) );
  AND2X4 U2152 ( .A(n2227), .B(n2026), .Y(n2226) );
  INVX4 U2153 ( .A(n2228), .Y(n2026) );
  AND2X4 U2154 ( .A(B[13]), .B(n2229), .Y(n2227) );
  OR2X4 U2155 ( .A(n131), .B(n2230), .Y(n2229) );
  OR2X4 U2156 ( .A(n2231), .B(n2232), .Y(n2230) );
  AND2X4 U2157 ( .A(n2233), .B(B[14]), .Y(n2232) );
  AND2X4 U2158 ( .A(A[2]), .B(n183), .Y(n2231) );
  AND2X4 U2159 ( .A(n2234), .B(n2228), .Y(n2225) );
  OR2X4 U2160 ( .A(n2235), .B(n2236), .Y(n2228) );
  OR2X4 U2161 ( .A(n2237), .B(n2238), .Y(n2236) );
  AND2X4 U2162 ( .A(B[14]), .B(n1210), .Y(n2238) );
  AND2X4 U2163 ( .A(n297), .B(A[0]), .Y(n2237) );
  AND2X4 U2164 ( .A(n183), .B(B[15]), .Y(n297) );
  OR2X4 U2165 ( .A(n2239), .B(n2240), .Y(n2235) );
  AND2X4 U2166 ( .A(n293), .B(A[1]), .Y(n2240) );
  AND2X4 U2167 ( .A(n182), .B(B[14]), .Y(n293) );
  INVX4 U2168 ( .A(B[15]), .Y(n182) );
  AND2X4 U2169 ( .A(n1207), .B(B[15]), .Y(n2239) );
  OR2X4 U2170 ( .A(n2241), .B(n2242), .Y(n2234) );
  OR2X4 U2171 ( .A(n137), .B(n2020), .Y(n2242) );
  OR2X4 U2172 ( .A(n2243), .B(n2244), .Y(n2241) );
  AND2X4 U2173 ( .A(n141), .B(B[14]), .Y(n2244) );
  AND2X4 U2174 ( .A(n142), .B(n183), .Y(n2243) );
  OR2X4 U2175 ( .A(n2245), .B(n2246), .Y(Y[14]) );
  AND2X4 U2176 ( .A(n2247), .B(n2248), .Y(n2246) );
  AND2X4 U2177 ( .A(n2249), .B(n2041), .Y(n2248) );
  OR2X4 U2178 ( .A(n2250), .B(n2251), .Y(n2041) );
  OR2X4 U2179 ( .A(n2252), .B(n2253), .Y(n2249) );
  INVX4 U2180 ( .A(n2040), .Y(n2247) );
  AND2X4 U2181 ( .A(n2040), .B(n2254), .Y(n2245) );
  OR2X4 U2182 ( .A(n2255), .B(n2039), .Y(n2254) );
  AND2X4 U2183 ( .A(n2251), .B(n2250), .Y(n2039) );
  AND2X4 U2184 ( .A(n2252), .B(n2253), .Y(n2255) );
  INVX4 U2185 ( .A(n2250), .Y(n2253) );
  AND2X4 U2186 ( .A(B[0]), .B(A[14]), .Y(n2250) );
  INVX4 U2187 ( .A(n2251), .Y(n2252) );
  OR2X4 U2188 ( .A(n2256), .B(n2257), .Y(n2251) );
  AND2X4 U2189 ( .A(n2258), .B(n2259), .Y(n2256) );
  OR2X4 U2190 ( .A(n2260), .B(n2261), .Y(n2040) );
  AND2X4 U2191 ( .A(n2262), .B(n2263), .Y(n2261) );
  AND2X4 U2192 ( .A(n2264), .B(n2056), .Y(n2263) );
  OR2X4 U2193 ( .A(n2265), .B(n2266), .Y(n2056) );
  OR2X4 U2194 ( .A(n2267), .B(n2268), .Y(n2264) );
  INVX4 U2195 ( .A(n2055), .Y(n2262) );
  AND2X4 U2196 ( .A(n2055), .B(n2269), .Y(n2260) );
  OR2X4 U2197 ( .A(n2270), .B(n2054), .Y(n2269) );
  AND2X4 U2198 ( .A(n2266), .B(n2265), .Y(n2054) );
  AND2X4 U2199 ( .A(n2267), .B(n2268), .Y(n2270) );
  INVX4 U2200 ( .A(n2265), .Y(n2268) );
  AND2X4 U2201 ( .A(B[1]), .B(A[13]), .Y(n2265) );
  INVX4 U2202 ( .A(n2266), .Y(n2267) );
  OR2X4 U2203 ( .A(n2271), .B(n2272), .Y(n2266) );
  AND2X4 U2204 ( .A(n2273), .B(n2274), .Y(n2271) );
  OR2X4 U2205 ( .A(n2275), .B(n2276), .Y(n2055) );
  AND2X4 U2206 ( .A(n2277), .B(n2278), .Y(n2276) );
  AND2X4 U2207 ( .A(n2279), .B(n2071), .Y(n2278) );
  OR2X4 U2208 ( .A(n2280), .B(n2281), .Y(n2071) );
  OR2X4 U2209 ( .A(n2282), .B(n2283), .Y(n2279) );
  INVX4 U2210 ( .A(n2070), .Y(n2277) );
  AND2X4 U2211 ( .A(n2070), .B(n2284), .Y(n2275) );
  OR2X4 U2212 ( .A(n2285), .B(n2069), .Y(n2284) );
  AND2X4 U2213 ( .A(n2281), .B(n2280), .Y(n2069) );
  AND2X4 U2214 ( .A(n2282), .B(n2283), .Y(n2285) );
  INVX4 U2215 ( .A(n2280), .Y(n2283) );
  AND2X4 U2216 ( .A(B[2]), .B(A[12]), .Y(n2280) );
  INVX4 U2217 ( .A(n2281), .Y(n2282) );
  OR2X4 U2218 ( .A(n2286), .B(n2287), .Y(n2281) );
  AND2X4 U2219 ( .A(n2288), .B(n2289), .Y(n2286) );
  OR2X4 U2220 ( .A(n2290), .B(n2291), .Y(n2070) );
  AND2X4 U2221 ( .A(n2292), .B(n2293), .Y(n2291) );
  AND2X4 U2222 ( .A(n2294), .B(n2086), .Y(n2293) );
  OR2X4 U2223 ( .A(n2295), .B(n2296), .Y(n2086) );
  OR2X4 U2224 ( .A(n2297), .B(n2298), .Y(n2294) );
  INVX4 U2225 ( .A(n2085), .Y(n2292) );
  AND2X4 U2226 ( .A(n2085), .B(n2299), .Y(n2290) );
  OR2X4 U2227 ( .A(n2300), .B(n2084), .Y(n2299) );
  AND2X4 U2228 ( .A(n2296), .B(n2295), .Y(n2084) );
  AND2X4 U2229 ( .A(n2297), .B(n2298), .Y(n2300) );
  INVX4 U2230 ( .A(n2295), .Y(n2298) );
  AND2X4 U2231 ( .A(B[3]), .B(A[11]), .Y(n2295) );
  INVX4 U2232 ( .A(n2296), .Y(n2297) );
  OR2X4 U2233 ( .A(n2301), .B(n2302), .Y(n2296) );
  AND2X4 U2234 ( .A(n2303), .B(n2304), .Y(n2301) );
  OR2X4 U2235 ( .A(n2305), .B(n2306), .Y(n2085) );
  AND2X4 U2236 ( .A(n2307), .B(n2308), .Y(n2306) );
  AND2X4 U2237 ( .A(n2309), .B(n2101), .Y(n2308) );
  OR2X4 U2238 ( .A(n2310), .B(n2311), .Y(n2101) );
  OR2X4 U2239 ( .A(n2312), .B(n2313), .Y(n2309) );
  INVX4 U2240 ( .A(n2100), .Y(n2307) );
  AND2X4 U2241 ( .A(n2100), .B(n2314), .Y(n2305) );
  OR2X4 U2242 ( .A(n2315), .B(n2099), .Y(n2314) );
  AND2X4 U2243 ( .A(n2311), .B(n2310), .Y(n2099) );
  AND2X4 U2244 ( .A(n2312), .B(n2313), .Y(n2315) );
  INVX4 U2245 ( .A(n2310), .Y(n2313) );
  AND2X4 U2246 ( .A(B[4]), .B(A[10]), .Y(n2310) );
  INVX4 U2247 ( .A(n2311), .Y(n2312) );
  OR2X4 U2248 ( .A(n2316), .B(n2317), .Y(n2311) );
  AND2X4 U2249 ( .A(n2318), .B(n2319), .Y(n2316) );
  OR2X4 U2250 ( .A(n2320), .B(n2321), .Y(n2100) );
  AND2X4 U2251 ( .A(n2322), .B(n2323), .Y(n2321) );
  AND2X4 U2252 ( .A(n2324), .B(n2116), .Y(n2323) );
  OR2X4 U2253 ( .A(n2325), .B(n2326), .Y(n2116) );
  OR2X4 U2254 ( .A(n2327), .B(n2328), .Y(n2324) );
  INVX4 U2255 ( .A(n2115), .Y(n2322) );
  AND2X4 U2256 ( .A(n2115), .B(n2329), .Y(n2320) );
  OR2X4 U2257 ( .A(n2330), .B(n2114), .Y(n2329) );
  AND2X4 U2258 ( .A(n2326), .B(n2325), .Y(n2114) );
  AND2X4 U2259 ( .A(n2327), .B(n2328), .Y(n2330) );
  INVX4 U2260 ( .A(n2325), .Y(n2328) );
  AND2X4 U2261 ( .A(B[5]), .B(A[9]), .Y(n2325) );
  INVX4 U2262 ( .A(n2326), .Y(n2327) );
  OR2X4 U2263 ( .A(n2331), .B(n2332), .Y(n2326) );
  AND2X4 U2264 ( .A(n2333), .B(n2334), .Y(n2331) );
  OR2X4 U2265 ( .A(n2335), .B(n2336), .Y(n2115) );
  AND2X4 U2266 ( .A(n2337), .B(n2338), .Y(n2336) );
  AND2X4 U2267 ( .A(n2339), .B(n2131), .Y(n2338) );
  OR2X4 U2268 ( .A(n2340), .B(n2341), .Y(n2131) );
  OR2X4 U2269 ( .A(n2342), .B(n2343), .Y(n2339) );
  INVX4 U2270 ( .A(n2130), .Y(n2337) );
  AND2X4 U2271 ( .A(n2130), .B(n2344), .Y(n2335) );
  OR2X4 U2272 ( .A(n2345), .B(n2129), .Y(n2344) );
  AND2X4 U2273 ( .A(n2341), .B(n2340), .Y(n2129) );
  AND2X4 U2274 ( .A(n2342), .B(n2343), .Y(n2345) );
  INVX4 U2275 ( .A(n2340), .Y(n2343) );
  AND2X4 U2276 ( .A(B[6]), .B(A[8]), .Y(n2340) );
  INVX4 U2277 ( .A(n2341), .Y(n2342) );
  OR2X4 U2278 ( .A(n2346), .B(n2347), .Y(n2341) );
  AND2X4 U2279 ( .A(n2348), .B(n2349), .Y(n2346) );
  OR2X4 U2280 ( .A(n2350), .B(n2351), .Y(n2130) );
  AND2X4 U2281 ( .A(n2352), .B(n2353), .Y(n2351) );
  AND2X4 U2282 ( .A(n2354), .B(n2146), .Y(n2353) );
  OR2X4 U2283 ( .A(n2355), .B(n2356), .Y(n2146) );
  OR2X4 U2284 ( .A(n2357), .B(n2358), .Y(n2354) );
  INVX4 U2285 ( .A(n2145), .Y(n2352) );
  AND2X4 U2286 ( .A(n2145), .B(n2359), .Y(n2350) );
  OR2X4 U2287 ( .A(n2360), .B(n2144), .Y(n2359) );
  AND2X4 U2288 ( .A(n2356), .B(n2355), .Y(n2144) );
  AND2X4 U2289 ( .A(n2357), .B(n2358), .Y(n2360) );
  INVX4 U2290 ( .A(n2355), .Y(n2358) );
  AND2X4 U2291 ( .A(B[7]), .B(A[7]), .Y(n2355) );
  INVX4 U2292 ( .A(n2356), .Y(n2357) );
  OR2X4 U2293 ( .A(n2361), .B(n2362), .Y(n2356) );
  AND2X4 U2294 ( .A(n2363), .B(n2364), .Y(n2361) );
  OR2X4 U2295 ( .A(n2365), .B(n2366), .Y(n2145) );
  AND2X4 U2296 ( .A(n2367), .B(n2368), .Y(n2366) );
  AND2X4 U2297 ( .A(n2369), .B(n2161), .Y(n2368) );
  OR2X4 U2298 ( .A(n2370), .B(n2371), .Y(n2161) );
  OR2X4 U2299 ( .A(n2372), .B(n2373), .Y(n2369) );
  INVX4 U2300 ( .A(n2160), .Y(n2367) );
  AND2X4 U2301 ( .A(n2160), .B(n2374), .Y(n2365) );
  OR2X4 U2302 ( .A(n2375), .B(n2159), .Y(n2374) );
  AND2X4 U2303 ( .A(n2371), .B(n2370), .Y(n2159) );
  AND2X4 U2304 ( .A(n2372), .B(n2373), .Y(n2375) );
  INVX4 U2305 ( .A(n2370), .Y(n2373) );
  AND2X4 U2306 ( .A(B[8]), .B(A[6]), .Y(n2370) );
  INVX4 U2307 ( .A(n2371), .Y(n2372) );
  OR2X4 U2308 ( .A(n2376), .B(n2377), .Y(n2371) );
  AND2X4 U2309 ( .A(n2378), .B(n2379), .Y(n2376) );
  OR2X4 U2310 ( .A(n2380), .B(n2381), .Y(n2160) );
  AND2X4 U2311 ( .A(n2382), .B(n2383), .Y(n2381) );
  AND2X4 U2312 ( .A(n2384), .B(n2176), .Y(n2383) );
  OR2X4 U2313 ( .A(n2385), .B(n2386), .Y(n2176) );
  OR2X4 U2314 ( .A(n2387), .B(n2388), .Y(n2384) );
  INVX4 U2315 ( .A(n2175), .Y(n2382) );
  AND2X4 U2316 ( .A(n2175), .B(n2389), .Y(n2380) );
  OR2X4 U2317 ( .A(n2390), .B(n2174), .Y(n2389) );
  AND2X4 U2318 ( .A(n2386), .B(n2385), .Y(n2174) );
  AND2X4 U2319 ( .A(n2387), .B(n2388), .Y(n2390) );
  INVX4 U2320 ( .A(n2385), .Y(n2388) );
  AND2X4 U2321 ( .A(B[9]), .B(A[5]), .Y(n2385) );
  INVX4 U2322 ( .A(n2386), .Y(n2387) );
  OR2X4 U2323 ( .A(n2391), .B(n2392), .Y(n2386) );
  AND2X4 U2324 ( .A(n2393), .B(n2394), .Y(n2391) );
  OR2X4 U2325 ( .A(n2395), .B(n2396), .Y(n2175) );
  AND2X4 U2326 ( .A(n2397), .B(n2398), .Y(n2396) );
  AND2X4 U2327 ( .A(n2399), .B(n2191), .Y(n2398) );
  OR2X4 U2328 ( .A(n2400), .B(n2401), .Y(n2191) );
  OR2X4 U2329 ( .A(n2402), .B(n2403), .Y(n2399) );
  INVX4 U2330 ( .A(n2190), .Y(n2397) );
  AND2X4 U2331 ( .A(n2190), .B(n2404), .Y(n2395) );
  OR2X4 U2332 ( .A(n2405), .B(n2189), .Y(n2404) );
  AND2X4 U2333 ( .A(n2401), .B(n2400), .Y(n2189) );
  AND2X4 U2334 ( .A(n2402), .B(n2403), .Y(n2405) );
  INVX4 U2335 ( .A(n2400), .Y(n2403) );
  AND2X4 U2336 ( .A(A[4]), .B(B[10]), .Y(n2400) );
  INVX4 U2337 ( .A(n2401), .Y(n2402) );
  OR2X4 U2338 ( .A(n2406), .B(n2407), .Y(n2401) );
  AND2X4 U2339 ( .A(n2408), .B(n2409), .Y(n2406) );
  OR2X4 U2340 ( .A(n2410), .B(n2411), .Y(n2409) );
  OR2X4 U2341 ( .A(n2412), .B(n2413), .Y(n2190) );
  AND2X4 U2342 ( .A(n2414), .B(n2415), .Y(n2413) );
  INVX4 U2343 ( .A(n2205), .Y(n2415) );
  OR2X4 U2344 ( .A(n2416), .B(n2417), .Y(n2414) );
  AND2X4 U2345 ( .A(n2207), .B(n2418), .Y(n2417) );
  AND2X4 U2346 ( .A(n2208), .B(n2419), .Y(n2416) );
  AND2X4 U2347 ( .A(n2205), .B(n2420), .Y(n2412) );
  OR2X4 U2348 ( .A(n2421), .B(n2204), .Y(n2420) );
  AND2X4 U2349 ( .A(n2207), .B(n2208), .Y(n2204) );
  INVX4 U2350 ( .A(n2418), .Y(n2208) );
  AND2X4 U2351 ( .A(n2419), .B(n2418), .Y(n2421) );
  OR2X4 U2352 ( .A(n2422), .B(n2423), .Y(n2418) );
  AND2X4 U2353 ( .A(n2424), .B(n2425), .Y(n2422) );
  OR2X4 U2354 ( .A(n2426), .B(n269), .Y(n2425) );
  AND2X4 U2355 ( .A(n2024), .B(n2427), .Y(n2426) );
  OR2X4 U2356 ( .A(n2428), .B(n1804), .Y(n2427) );
  OR2X4 U2357 ( .A(n2428), .B(n142), .Y(n2424) );
  INVX4 U2358 ( .A(n2207), .Y(n2419) );
  AND2X4 U2359 ( .A(A[3]), .B(B[11]), .Y(n2207) );
  OR2X4 U2360 ( .A(n2429), .B(n2430), .Y(n2205) );
  AND2X4 U2361 ( .A(n2431), .B(n2224), .Y(n2430) );
  INVX4 U2362 ( .A(n2432), .Y(n2224) );
  AND2X4 U2363 ( .A(B[12]), .B(n2433), .Y(n2431) );
  OR2X4 U2364 ( .A(n131), .B(n2434), .Y(n2433) );
  OR2X4 U2365 ( .A(n2435), .B(n2436), .Y(n2434) );
  AND2X4 U2366 ( .A(n2233), .B(B[13]), .Y(n2436) );
  AND2X4 U2367 ( .A(A[2]), .B(n2020), .Y(n2435) );
  AND2X4 U2368 ( .A(n2437), .B(n2432), .Y(n2429) );
  OR2X4 U2369 ( .A(n2438), .B(n2439), .Y(n2432) );
  AND2X4 U2370 ( .A(B[14]), .B(n2440), .Y(n2439) );
  OR2X4 U2371 ( .A(n2441), .B(n1207), .Y(n2440) );
  AND2X4 U2372 ( .A(A[0]), .B(n2020), .Y(n2441) );
  AND2X4 U2373 ( .A(B[13]), .B(n2442), .Y(n2438) );
  OR2X4 U2374 ( .A(n2443), .B(n1210), .Y(n2442) );
  AND2X4 U2375 ( .A(A[1]), .B(n183), .Y(n2443) );
  INVX4 U2376 ( .A(B[14]), .Y(n183) );
  OR2X4 U2377 ( .A(n2444), .B(n2445), .Y(n2437) );
  OR2X4 U2378 ( .A(n137), .B(n269), .Y(n2445) );
  OR2X4 U2379 ( .A(n2446), .B(n2447), .Y(n2444) );
  AND2X4 U2380 ( .A(n141), .B(B[13]), .Y(n2447) );
  AND2X4 U2381 ( .A(n142), .B(n2020), .Y(n2446) );
  OR2X4 U2382 ( .A(n2448), .B(n2449), .Y(Y[13]) );
  AND2X4 U2383 ( .A(n2450), .B(n2451), .Y(n2449) );
  AND2X4 U2384 ( .A(n2452), .B(n2259), .Y(n2451) );
  OR2X4 U2385 ( .A(n2453), .B(n2454), .Y(n2259) );
  OR2X4 U2386 ( .A(n2455), .B(n2456), .Y(n2452) );
  INVX4 U2387 ( .A(n2258), .Y(n2450) );
  AND2X4 U2388 ( .A(n2258), .B(n2457), .Y(n2448) );
  OR2X4 U2389 ( .A(n2458), .B(n2257), .Y(n2457) );
  AND2X4 U2390 ( .A(n2454), .B(n2453), .Y(n2257) );
  AND2X4 U2391 ( .A(n2455), .B(n2456), .Y(n2458) );
  INVX4 U2392 ( .A(n2453), .Y(n2456) );
  AND2X4 U2393 ( .A(B[0]), .B(A[13]), .Y(n2453) );
  INVX4 U2394 ( .A(n2454), .Y(n2455) );
  OR2X4 U2395 ( .A(n2459), .B(n2460), .Y(n2454) );
  AND2X4 U2396 ( .A(n2461), .B(n2462), .Y(n2459) );
  OR2X4 U2397 ( .A(n2463), .B(n2464), .Y(n2258) );
  AND2X4 U2398 ( .A(n2465), .B(n2466), .Y(n2464) );
  AND2X4 U2399 ( .A(n2467), .B(n2274), .Y(n2466) );
  OR2X4 U2400 ( .A(n2468), .B(n2469), .Y(n2274) );
  OR2X4 U2401 ( .A(n2470), .B(n2471), .Y(n2467) );
  INVX4 U2402 ( .A(n2273), .Y(n2465) );
  AND2X4 U2403 ( .A(n2273), .B(n2472), .Y(n2463) );
  OR2X4 U2404 ( .A(n2473), .B(n2272), .Y(n2472) );
  AND2X4 U2405 ( .A(n2469), .B(n2468), .Y(n2272) );
  AND2X4 U2406 ( .A(n2470), .B(n2471), .Y(n2473) );
  INVX4 U2407 ( .A(n2468), .Y(n2471) );
  AND2X4 U2408 ( .A(B[1]), .B(A[12]), .Y(n2468) );
  INVX4 U2409 ( .A(n2469), .Y(n2470) );
  OR2X4 U2410 ( .A(n2474), .B(n2475), .Y(n2469) );
  AND2X4 U2411 ( .A(n2476), .B(n2477), .Y(n2474) );
  OR2X4 U2412 ( .A(n2478), .B(n2479), .Y(n2273) );
  AND2X4 U2413 ( .A(n2480), .B(n2481), .Y(n2479) );
  AND2X4 U2414 ( .A(n2482), .B(n2289), .Y(n2481) );
  OR2X4 U2415 ( .A(n2483), .B(n2484), .Y(n2289) );
  OR2X4 U2416 ( .A(n2485), .B(n2486), .Y(n2482) );
  INVX4 U2417 ( .A(n2288), .Y(n2480) );
  AND2X4 U2418 ( .A(n2288), .B(n2487), .Y(n2478) );
  OR2X4 U2419 ( .A(n2488), .B(n2287), .Y(n2487) );
  AND2X4 U2420 ( .A(n2484), .B(n2483), .Y(n2287) );
  AND2X4 U2421 ( .A(n2485), .B(n2486), .Y(n2488) );
  INVX4 U2422 ( .A(n2483), .Y(n2486) );
  AND2X4 U2423 ( .A(B[2]), .B(A[11]), .Y(n2483) );
  INVX4 U2424 ( .A(n2484), .Y(n2485) );
  OR2X4 U2425 ( .A(n2489), .B(n2490), .Y(n2484) );
  AND2X4 U2426 ( .A(n2491), .B(n2492), .Y(n2489) );
  OR2X4 U2427 ( .A(n2493), .B(n2494), .Y(n2288) );
  AND2X4 U2428 ( .A(n2495), .B(n2496), .Y(n2494) );
  AND2X4 U2429 ( .A(n2497), .B(n2304), .Y(n2496) );
  OR2X4 U2430 ( .A(n2498), .B(n2499), .Y(n2304) );
  OR2X4 U2431 ( .A(n2500), .B(n2501), .Y(n2497) );
  INVX4 U2432 ( .A(n2303), .Y(n2495) );
  AND2X4 U2433 ( .A(n2303), .B(n2502), .Y(n2493) );
  OR2X4 U2434 ( .A(n2503), .B(n2302), .Y(n2502) );
  AND2X4 U2435 ( .A(n2499), .B(n2498), .Y(n2302) );
  AND2X4 U2436 ( .A(n2500), .B(n2501), .Y(n2503) );
  INVX4 U2437 ( .A(n2498), .Y(n2501) );
  AND2X4 U2438 ( .A(B[3]), .B(A[10]), .Y(n2498) );
  INVX4 U2439 ( .A(n2499), .Y(n2500) );
  OR2X4 U2440 ( .A(n2504), .B(n2505), .Y(n2499) );
  AND2X4 U2441 ( .A(n2506), .B(n2507), .Y(n2504) );
  OR2X4 U2442 ( .A(n2508), .B(n2509), .Y(n2303) );
  AND2X4 U2443 ( .A(n2510), .B(n2511), .Y(n2509) );
  AND2X4 U2444 ( .A(n2512), .B(n2319), .Y(n2511) );
  OR2X4 U2445 ( .A(n2513), .B(n2514), .Y(n2319) );
  OR2X4 U2446 ( .A(n2515), .B(n2516), .Y(n2512) );
  INVX4 U2447 ( .A(n2318), .Y(n2510) );
  AND2X4 U2448 ( .A(n2318), .B(n2517), .Y(n2508) );
  OR2X4 U2449 ( .A(n2518), .B(n2317), .Y(n2517) );
  AND2X4 U2450 ( .A(n2514), .B(n2513), .Y(n2317) );
  AND2X4 U2451 ( .A(n2515), .B(n2516), .Y(n2518) );
  INVX4 U2452 ( .A(n2513), .Y(n2516) );
  AND2X4 U2453 ( .A(B[4]), .B(A[9]), .Y(n2513) );
  INVX4 U2454 ( .A(n2514), .Y(n2515) );
  OR2X4 U2455 ( .A(n2519), .B(n2520), .Y(n2514) );
  AND2X4 U2456 ( .A(n2521), .B(n2522), .Y(n2519) );
  OR2X4 U2457 ( .A(n2523), .B(n2524), .Y(n2318) );
  AND2X4 U2458 ( .A(n2525), .B(n2526), .Y(n2524) );
  AND2X4 U2459 ( .A(n2527), .B(n2334), .Y(n2526) );
  OR2X4 U2460 ( .A(n2528), .B(n2529), .Y(n2334) );
  OR2X4 U2461 ( .A(n2530), .B(n2531), .Y(n2527) );
  INVX4 U2462 ( .A(n2333), .Y(n2525) );
  AND2X4 U2463 ( .A(n2333), .B(n2532), .Y(n2523) );
  OR2X4 U2464 ( .A(n2533), .B(n2332), .Y(n2532) );
  AND2X4 U2465 ( .A(n2529), .B(n2528), .Y(n2332) );
  AND2X4 U2466 ( .A(n2530), .B(n2531), .Y(n2533) );
  INVX4 U2467 ( .A(n2528), .Y(n2531) );
  AND2X4 U2468 ( .A(B[5]), .B(A[8]), .Y(n2528) );
  INVX4 U2469 ( .A(n2529), .Y(n2530) );
  OR2X4 U2470 ( .A(n2534), .B(n2535), .Y(n2529) );
  AND2X4 U2471 ( .A(n2536), .B(n2537), .Y(n2534) );
  OR2X4 U2472 ( .A(n2538), .B(n2539), .Y(n2333) );
  AND2X4 U2473 ( .A(n2540), .B(n2541), .Y(n2539) );
  AND2X4 U2474 ( .A(n2542), .B(n2349), .Y(n2541) );
  OR2X4 U2475 ( .A(n2543), .B(n2544), .Y(n2349) );
  OR2X4 U2476 ( .A(n2545), .B(n2546), .Y(n2542) );
  INVX4 U2477 ( .A(n2348), .Y(n2540) );
  AND2X4 U2478 ( .A(n2348), .B(n2547), .Y(n2538) );
  OR2X4 U2479 ( .A(n2548), .B(n2347), .Y(n2547) );
  AND2X4 U2480 ( .A(n2544), .B(n2543), .Y(n2347) );
  AND2X4 U2481 ( .A(n2545), .B(n2546), .Y(n2548) );
  INVX4 U2482 ( .A(n2543), .Y(n2546) );
  AND2X4 U2483 ( .A(B[6]), .B(A[7]), .Y(n2543) );
  INVX4 U2484 ( .A(n2544), .Y(n2545) );
  OR2X4 U2485 ( .A(n2549), .B(n2550), .Y(n2544) );
  AND2X4 U2486 ( .A(n2551), .B(n2552), .Y(n2549) );
  OR2X4 U2487 ( .A(n2553), .B(n2554), .Y(n2348) );
  AND2X4 U2488 ( .A(n2555), .B(n2556), .Y(n2554) );
  AND2X4 U2489 ( .A(n2557), .B(n2364), .Y(n2556) );
  OR2X4 U2490 ( .A(n2558), .B(n2559), .Y(n2364) );
  OR2X4 U2491 ( .A(n2560), .B(n2561), .Y(n2557) );
  INVX4 U2492 ( .A(n2363), .Y(n2555) );
  AND2X4 U2493 ( .A(n2363), .B(n2562), .Y(n2553) );
  OR2X4 U2494 ( .A(n2563), .B(n2362), .Y(n2562) );
  AND2X4 U2495 ( .A(n2559), .B(n2558), .Y(n2362) );
  AND2X4 U2496 ( .A(n2560), .B(n2561), .Y(n2563) );
  INVX4 U2497 ( .A(n2558), .Y(n2561) );
  AND2X4 U2498 ( .A(B[7]), .B(A[6]), .Y(n2558) );
  INVX4 U2499 ( .A(n2559), .Y(n2560) );
  OR2X4 U2500 ( .A(n2564), .B(n2565), .Y(n2559) );
  AND2X4 U2501 ( .A(n2566), .B(n2567), .Y(n2564) );
  OR2X4 U2502 ( .A(n2568), .B(n2569), .Y(n2363) );
  AND2X4 U2503 ( .A(n2570), .B(n2571), .Y(n2569) );
  AND2X4 U2504 ( .A(n2572), .B(n2379), .Y(n2571) );
  OR2X4 U2505 ( .A(n2573), .B(n2574), .Y(n2379) );
  OR2X4 U2506 ( .A(n2575), .B(n2576), .Y(n2572) );
  INVX4 U2507 ( .A(n2378), .Y(n2570) );
  AND2X4 U2508 ( .A(n2378), .B(n2577), .Y(n2568) );
  OR2X4 U2509 ( .A(n2578), .B(n2377), .Y(n2577) );
  AND2X4 U2510 ( .A(n2574), .B(n2573), .Y(n2377) );
  AND2X4 U2511 ( .A(n2575), .B(n2576), .Y(n2578) );
  INVX4 U2512 ( .A(n2573), .Y(n2576) );
  AND2X4 U2513 ( .A(B[8]), .B(A[5]), .Y(n2573) );
  INVX4 U2514 ( .A(n2574), .Y(n2575) );
  OR2X4 U2515 ( .A(n2579), .B(n2580), .Y(n2574) );
  AND2X4 U2516 ( .A(n2581), .B(n2582), .Y(n2579) );
  OR2X4 U2517 ( .A(n2583), .B(n2584), .Y(n2378) );
  AND2X4 U2518 ( .A(n2585), .B(n2586), .Y(n2584) );
  AND2X4 U2519 ( .A(n2587), .B(n2394), .Y(n2586) );
  OR2X4 U2520 ( .A(n2588), .B(n2589), .Y(n2394) );
  OR2X4 U2521 ( .A(n2590), .B(n2591), .Y(n2587) );
  INVX4 U2522 ( .A(n2393), .Y(n2585) );
  AND2X4 U2523 ( .A(n2393), .B(n2592), .Y(n2583) );
  OR2X4 U2524 ( .A(n2593), .B(n2392), .Y(n2592) );
  AND2X4 U2525 ( .A(n2589), .B(n2588), .Y(n2392) );
  AND2X4 U2526 ( .A(n2590), .B(n2591), .Y(n2593) );
  INVX4 U2527 ( .A(n2588), .Y(n2591) );
  AND2X4 U2528 ( .A(B[9]), .B(A[4]), .Y(n2588) );
  INVX4 U2529 ( .A(n2589), .Y(n2590) );
  OR2X4 U2530 ( .A(n2594), .B(n2595), .Y(n2589) );
  AND2X4 U2531 ( .A(n2596), .B(n2597), .Y(n2594) );
  OR2X4 U2532 ( .A(n2598), .B(n2599), .Y(n2597) );
  OR2X4 U2533 ( .A(n2600), .B(n2601), .Y(n2393) );
  AND2X4 U2534 ( .A(n2602), .B(n2603), .Y(n2601) );
  INVX4 U2535 ( .A(n2408), .Y(n2603) );
  OR2X4 U2536 ( .A(n2604), .B(n2605), .Y(n2602) );
  AND2X4 U2537 ( .A(n2410), .B(n2606), .Y(n2605) );
  AND2X4 U2538 ( .A(n2411), .B(n2607), .Y(n2604) );
  AND2X4 U2539 ( .A(n2408), .B(n2608), .Y(n2600) );
  OR2X4 U2540 ( .A(n2609), .B(n2407), .Y(n2608) );
  AND2X4 U2541 ( .A(n2410), .B(n2411), .Y(n2407) );
  INVX4 U2542 ( .A(n2606), .Y(n2411) );
  AND2X4 U2543 ( .A(n2607), .B(n2606), .Y(n2609) );
  OR2X4 U2544 ( .A(n2610), .B(n423), .Y(n2606) );
  AND2X4 U2545 ( .A(n2611), .B(n2612), .Y(n2610) );
  OR2X4 U2546 ( .A(n2613), .B(n2423), .Y(n2612) );
  AND2X4 U2547 ( .A(n2024), .B(n2614), .Y(n2613) );
  OR2X4 U2548 ( .A(n2615), .B(n1804), .Y(n2614) );
  OR2X4 U2549 ( .A(n2615), .B(n142), .Y(n2611) );
  INVX4 U2550 ( .A(n2410), .Y(n2607) );
  AND2X4 U2551 ( .A(A[3]), .B(B[10]), .Y(n2410) );
  OR2X4 U2552 ( .A(n2616), .B(n2617), .Y(n2408) );
  AND2X4 U2553 ( .A(n2618), .B(n2428), .Y(n2617) );
  INVX4 U2554 ( .A(n2619), .Y(n2428) );
  AND2X4 U2555 ( .A(B[11]), .B(n2620), .Y(n2618) );
  OR2X4 U2556 ( .A(n131), .B(n2621), .Y(n2620) );
  OR2X4 U2557 ( .A(n2622), .B(n2623), .Y(n2621) );
  AND2X4 U2558 ( .A(n2233), .B(B[12]), .Y(n2623) );
  AND2X4 U2559 ( .A(A[2]), .B(n269), .Y(n2622) );
  AND2X4 U2560 ( .A(n2624), .B(n2619), .Y(n2616) );
  OR2X4 U2561 ( .A(n2625), .B(n2626), .Y(n2619) );
  AND2X4 U2562 ( .A(B[13]), .B(n2627), .Y(n2626) );
  OR2X4 U2563 ( .A(n2628), .B(n1207), .Y(n2627) );
  AND2X4 U2564 ( .A(A[0]), .B(n269), .Y(n2628) );
  AND2X4 U2565 ( .A(B[12]), .B(n2629), .Y(n2625) );
  OR2X4 U2566 ( .A(n2630), .B(n1210), .Y(n2629) );
  AND2X4 U2567 ( .A(A[1]), .B(n2020), .Y(n2630) );
  INVX4 U2568 ( .A(B[13]), .Y(n2020) );
  OR2X4 U2569 ( .A(n2631), .B(n2632), .Y(n2624) );
  OR2X4 U2570 ( .A(n137), .B(n2423), .Y(n2632) );
  OR2X4 U2571 ( .A(n2633), .B(n2634), .Y(n2631) );
  AND2X4 U2572 ( .A(n141), .B(B[12]), .Y(n2634) );
  AND2X4 U2573 ( .A(n142), .B(n269), .Y(n2633) );
  OR2X4 U2574 ( .A(n2635), .B(n2636), .Y(Y[12]) );
  AND2X4 U2575 ( .A(n2637), .B(n2638), .Y(n2636) );
  AND2X4 U2576 ( .A(n2639), .B(n2462), .Y(n2638) );
  OR2X4 U2577 ( .A(n2640), .B(n2641), .Y(n2462) );
  OR2X4 U2578 ( .A(n2642), .B(n2643), .Y(n2639) );
  INVX4 U2579 ( .A(n2461), .Y(n2637) );
  AND2X4 U2580 ( .A(n2461), .B(n2644), .Y(n2635) );
  OR2X4 U2581 ( .A(n2645), .B(n2460), .Y(n2644) );
  AND2X4 U2582 ( .A(n2641), .B(n2640), .Y(n2460) );
  AND2X4 U2583 ( .A(n2642), .B(n2643), .Y(n2645) );
  INVX4 U2584 ( .A(n2640), .Y(n2643) );
  AND2X4 U2585 ( .A(B[0]), .B(A[12]), .Y(n2640) );
  INVX4 U2586 ( .A(n2641), .Y(n2642) );
  OR2X4 U2587 ( .A(n2646), .B(n2647), .Y(n2641) );
  AND2X4 U2588 ( .A(n2648), .B(n2649), .Y(n2646) );
  OR2X4 U2589 ( .A(n2650), .B(n2651), .Y(n2461) );
  AND2X4 U2590 ( .A(n2652), .B(n2653), .Y(n2651) );
  AND2X4 U2591 ( .A(n2654), .B(n2477), .Y(n2653) );
  OR2X4 U2592 ( .A(n2655), .B(n2656), .Y(n2477) );
  OR2X4 U2593 ( .A(n2657), .B(n2658), .Y(n2654) );
  INVX4 U2594 ( .A(n2476), .Y(n2652) );
  AND2X4 U2595 ( .A(n2476), .B(n2659), .Y(n2650) );
  OR2X4 U2596 ( .A(n2660), .B(n2475), .Y(n2659) );
  AND2X4 U2597 ( .A(n2656), .B(n2655), .Y(n2475) );
  AND2X4 U2598 ( .A(n2657), .B(n2658), .Y(n2660) );
  INVX4 U2599 ( .A(n2655), .Y(n2658) );
  AND2X4 U2600 ( .A(B[1]), .B(A[11]), .Y(n2655) );
  INVX4 U2601 ( .A(n2656), .Y(n2657) );
  OR2X4 U2602 ( .A(n2661), .B(n2662), .Y(n2656) );
  AND2X4 U2603 ( .A(n2663), .B(n2664), .Y(n2661) );
  OR2X4 U2604 ( .A(n2665), .B(n2666), .Y(n2476) );
  AND2X4 U2605 ( .A(n2667), .B(n2668), .Y(n2666) );
  AND2X4 U2606 ( .A(n2669), .B(n2492), .Y(n2668) );
  OR2X4 U2607 ( .A(n2670), .B(n2671), .Y(n2492) );
  OR2X4 U2608 ( .A(n2672), .B(n2673), .Y(n2669) );
  INVX4 U2609 ( .A(n2491), .Y(n2667) );
  AND2X4 U2610 ( .A(n2491), .B(n2674), .Y(n2665) );
  OR2X4 U2611 ( .A(n2675), .B(n2490), .Y(n2674) );
  AND2X4 U2612 ( .A(n2671), .B(n2670), .Y(n2490) );
  AND2X4 U2613 ( .A(n2672), .B(n2673), .Y(n2675) );
  INVX4 U2614 ( .A(n2670), .Y(n2673) );
  AND2X4 U2615 ( .A(B[2]), .B(A[10]), .Y(n2670) );
  INVX4 U2616 ( .A(n2671), .Y(n2672) );
  OR2X4 U2617 ( .A(n2676), .B(n2677), .Y(n2671) );
  AND2X4 U2618 ( .A(n2678), .B(n2679), .Y(n2676) );
  OR2X4 U2619 ( .A(n2680), .B(n2681), .Y(n2491) );
  AND2X4 U2620 ( .A(n2682), .B(n2683), .Y(n2681) );
  AND2X4 U2621 ( .A(n2684), .B(n2507), .Y(n2683) );
  OR2X4 U2622 ( .A(n2685), .B(n2686), .Y(n2507) );
  OR2X4 U2623 ( .A(n2687), .B(n2688), .Y(n2684) );
  INVX4 U2624 ( .A(n2506), .Y(n2682) );
  AND2X4 U2625 ( .A(n2506), .B(n2689), .Y(n2680) );
  OR2X4 U2626 ( .A(n2690), .B(n2505), .Y(n2689) );
  AND2X4 U2627 ( .A(n2686), .B(n2685), .Y(n2505) );
  AND2X4 U2628 ( .A(n2687), .B(n2688), .Y(n2690) );
  INVX4 U2629 ( .A(n2685), .Y(n2688) );
  AND2X4 U2630 ( .A(B[3]), .B(A[9]), .Y(n2685) );
  INVX4 U2631 ( .A(n2686), .Y(n2687) );
  OR2X4 U2632 ( .A(n2691), .B(n2692), .Y(n2686) );
  AND2X4 U2633 ( .A(n2693), .B(n2694), .Y(n2691) );
  OR2X4 U2634 ( .A(n2695), .B(n2696), .Y(n2506) );
  AND2X4 U2635 ( .A(n2697), .B(n2698), .Y(n2696) );
  AND2X4 U2636 ( .A(n2699), .B(n2522), .Y(n2698) );
  OR2X4 U2637 ( .A(n2700), .B(n2701), .Y(n2522) );
  OR2X4 U2638 ( .A(n2702), .B(n2703), .Y(n2699) );
  INVX4 U2639 ( .A(n2521), .Y(n2697) );
  AND2X4 U2640 ( .A(n2521), .B(n2704), .Y(n2695) );
  OR2X4 U2641 ( .A(n2705), .B(n2520), .Y(n2704) );
  AND2X4 U2642 ( .A(n2701), .B(n2700), .Y(n2520) );
  AND2X4 U2643 ( .A(n2702), .B(n2703), .Y(n2705) );
  INVX4 U2644 ( .A(n2700), .Y(n2703) );
  AND2X4 U2645 ( .A(B[4]), .B(A[8]), .Y(n2700) );
  INVX4 U2646 ( .A(n2701), .Y(n2702) );
  OR2X4 U2647 ( .A(n2706), .B(n2707), .Y(n2701) );
  AND2X4 U2648 ( .A(n2708), .B(n2709), .Y(n2706) );
  OR2X4 U2649 ( .A(n2710), .B(n2711), .Y(n2521) );
  AND2X4 U2650 ( .A(n2712), .B(n2713), .Y(n2711) );
  AND2X4 U2651 ( .A(n2714), .B(n2537), .Y(n2713) );
  OR2X4 U2652 ( .A(n2715), .B(n2716), .Y(n2537) );
  OR2X4 U2653 ( .A(n2717), .B(n2718), .Y(n2714) );
  INVX4 U2654 ( .A(n2536), .Y(n2712) );
  AND2X4 U2655 ( .A(n2536), .B(n2719), .Y(n2710) );
  OR2X4 U2656 ( .A(n2720), .B(n2535), .Y(n2719) );
  AND2X4 U2657 ( .A(n2716), .B(n2715), .Y(n2535) );
  AND2X4 U2658 ( .A(n2717), .B(n2718), .Y(n2720) );
  INVX4 U2659 ( .A(n2715), .Y(n2718) );
  AND2X4 U2660 ( .A(B[5]), .B(A[7]), .Y(n2715) );
  INVX4 U2661 ( .A(n2716), .Y(n2717) );
  OR2X4 U2662 ( .A(n2721), .B(n2722), .Y(n2716) );
  AND2X4 U2663 ( .A(n2723), .B(n2724), .Y(n2721) );
  OR2X4 U2664 ( .A(n2725), .B(n2726), .Y(n2536) );
  AND2X4 U2665 ( .A(n2727), .B(n2728), .Y(n2726) );
  AND2X4 U2666 ( .A(n2729), .B(n2552), .Y(n2728) );
  OR2X4 U2667 ( .A(n2730), .B(n2731), .Y(n2552) );
  OR2X4 U2668 ( .A(n2732), .B(n2733), .Y(n2729) );
  INVX4 U2669 ( .A(n2551), .Y(n2727) );
  AND2X4 U2670 ( .A(n2551), .B(n2734), .Y(n2725) );
  OR2X4 U2671 ( .A(n2735), .B(n2550), .Y(n2734) );
  AND2X4 U2672 ( .A(n2731), .B(n2730), .Y(n2550) );
  AND2X4 U2673 ( .A(n2732), .B(n2733), .Y(n2735) );
  INVX4 U2674 ( .A(n2730), .Y(n2733) );
  AND2X4 U2675 ( .A(B[6]), .B(A[6]), .Y(n2730) );
  INVX4 U2676 ( .A(n2731), .Y(n2732) );
  OR2X4 U2677 ( .A(n2736), .B(n2737), .Y(n2731) );
  AND2X4 U2678 ( .A(n2738), .B(n2739), .Y(n2736) );
  OR2X4 U2679 ( .A(n2740), .B(n2741), .Y(n2551) );
  AND2X4 U2680 ( .A(n2742), .B(n2743), .Y(n2741) );
  AND2X4 U2681 ( .A(n2744), .B(n2567), .Y(n2743) );
  OR2X4 U2682 ( .A(n2745), .B(n2746), .Y(n2567) );
  OR2X4 U2683 ( .A(n2747), .B(n2748), .Y(n2744) );
  INVX4 U2684 ( .A(n2566), .Y(n2742) );
  AND2X4 U2685 ( .A(n2566), .B(n2749), .Y(n2740) );
  OR2X4 U2686 ( .A(n2750), .B(n2565), .Y(n2749) );
  AND2X4 U2687 ( .A(n2746), .B(n2745), .Y(n2565) );
  AND2X4 U2688 ( .A(n2747), .B(n2748), .Y(n2750) );
  INVX4 U2689 ( .A(n2745), .Y(n2748) );
  AND2X4 U2690 ( .A(B[7]), .B(A[5]), .Y(n2745) );
  INVX4 U2691 ( .A(n2746), .Y(n2747) );
  OR2X4 U2692 ( .A(n2751), .B(n2752), .Y(n2746) );
  AND2X4 U2693 ( .A(n2753), .B(n2754), .Y(n2751) );
  OR2X4 U2694 ( .A(n2755), .B(n2756), .Y(n2566) );
  AND2X4 U2695 ( .A(n2757), .B(n2758), .Y(n2756) );
  AND2X4 U2696 ( .A(n2759), .B(n2582), .Y(n2758) );
  OR2X4 U2697 ( .A(n2760), .B(n2761), .Y(n2582) );
  OR2X4 U2698 ( .A(n2762), .B(n2763), .Y(n2759) );
  INVX4 U2699 ( .A(n2581), .Y(n2757) );
  AND2X4 U2700 ( .A(n2581), .B(n2764), .Y(n2755) );
  OR2X4 U2701 ( .A(n2765), .B(n2580), .Y(n2764) );
  AND2X4 U2702 ( .A(n2761), .B(n2760), .Y(n2580) );
  AND2X4 U2703 ( .A(n2762), .B(n2763), .Y(n2765) );
  INVX4 U2704 ( .A(n2760), .Y(n2763) );
  AND2X4 U2705 ( .A(B[8]), .B(A[4]), .Y(n2760) );
  INVX4 U2706 ( .A(n2761), .Y(n2762) );
  OR2X4 U2707 ( .A(n2766), .B(n2767), .Y(n2761) );
  AND2X4 U2708 ( .A(n2768), .B(n2769), .Y(n2766) );
  OR2X4 U2709 ( .A(n2770), .B(n2771), .Y(n2769) );
  OR2X4 U2710 ( .A(n2772), .B(n2773), .Y(n2581) );
  AND2X4 U2711 ( .A(n2774), .B(n2775), .Y(n2773) );
  INVX4 U2712 ( .A(n2596), .Y(n2775) );
  OR2X4 U2713 ( .A(n2776), .B(n2777), .Y(n2774) );
  AND2X4 U2714 ( .A(n2598), .B(n2778), .Y(n2777) );
  AND2X4 U2715 ( .A(n2599), .B(n2779), .Y(n2776) );
  AND2X4 U2716 ( .A(n2596), .B(n2780), .Y(n2772) );
  OR2X4 U2717 ( .A(n2781), .B(n2595), .Y(n2780) );
  AND2X4 U2718 ( .A(n2598), .B(n2599), .Y(n2595) );
  INVX4 U2719 ( .A(n2778), .Y(n2599) );
  AND2X4 U2720 ( .A(n2779), .B(n2778), .Y(n2781) );
  OR2X4 U2721 ( .A(n2782), .B(n2783), .Y(n2778) );
  AND2X4 U2722 ( .A(n2784), .B(n2785), .Y(n2782) );
  OR2X4 U2723 ( .A(n2786), .B(n423), .Y(n2785) );
  AND2X4 U2724 ( .A(n2024), .B(n2787), .Y(n2786) );
  OR2X4 U2725 ( .A(n2788), .B(n1804), .Y(n2787) );
  OR2X4 U2726 ( .A(n2788), .B(n142), .Y(n2784) );
  INVX4 U2727 ( .A(n2598), .Y(n2779) );
  AND2X4 U2728 ( .A(A[3]), .B(B[9]), .Y(n2598) );
  OR2X4 U2729 ( .A(n2789), .B(n2790), .Y(n2596) );
  AND2X4 U2730 ( .A(n2791), .B(n2615), .Y(n2790) );
  INVX4 U2731 ( .A(n2792), .Y(n2615) );
  AND2X4 U2732 ( .A(B[10]), .B(n2793), .Y(n2791) );
  OR2X4 U2733 ( .A(n131), .B(n2794), .Y(n2793) );
  OR2X4 U2734 ( .A(n2795), .B(n2796), .Y(n2794) );
  AND2X4 U2735 ( .A(n2233), .B(B[11]), .Y(n2796) );
  AND2X4 U2736 ( .A(A[2]), .B(n2423), .Y(n2795) );
  AND2X4 U2737 ( .A(n2797), .B(n2792), .Y(n2789) );
  OR2X4 U2738 ( .A(n2798), .B(n2799), .Y(n2792) );
  AND2X4 U2739 ( .A(B[12]), .B(n2800), .Y(n2799) );
  OR2X4 U2740 ( .A(n2801), .B(n1207), .Y(n2800) );
  AND2X4 U2741 ( .A(A[0]), .B(n2423), .Y(n2801) );
  AND2X4 U2742 ( .A(B[11]), .B(n2802), .Y(n2798) );
  OR2X4 U2743 ( .A(n2803), .B(n1210), .Y(n2802) );
  AND2X4 U2744 ( .A(A[1]), .B(n269), .Y(n2803) );
  INVX4 U2745 ( .A(B[12]), .Y(n269) );
  OR2X4 U2746 ( .A(n2804), .B(n2805), .Y(n2797) );
  OR2X4 U2747 ( .A(n137), .B(n423), .Y(n2805) );
  OR2X4 U2748 ( .A(n2806), .B(n2807), .Y(n2804) );
  AND2X4 U2749 ( .A(n141), .B(B[11]), .Y(n2807) );
  AND2X4 U2750 ( .A(n142), .B(n2423), .Y(n2806) );
  OR2X4 U2751 ( .A(n2808), .B(n2809), .Y(Y[11]) );
  AND2X4 U2752 ( .A(n2810), .B(n2811), .Y(n2809) );
  AND2X4 U2753 ( .A(n2812), .B(n2649), .Y(n2811) );
  OR2X4 U2754 ( .A(n2813), .B(n2814), .Y(n2649) );
  OR2X4 U2755 ( .A(n2815), .B(n2816), .Y(n2812) );
  INVX4 U2756 ( .A(n2648), .Y(n2810) );
  AND2X4 U2757 ( .A(n2648), .B(n2817), .Y(n2808) );
  OR2X4 U2758 ( .A(n2818), .B(n2647), .Y(n2817) );
  AND2X4 U2759 ( .A(n2814), .B(n2813), .Y(n2647) );
  AND2X4 U2760 ( .A(n2815), .B(n2816), .Y(n2818) );
  INVX4 U2761 ( .A(n2813), .Y(n2816) );
  AND2X4 U2762 ( .A(B[0]), .B(A[11]), .Y(n2813) );
  INVX4 U2763 ( .A(n2814), .Y(n2815) );
  OR2X4 U2764 ( .A(n2819), .B(n2820), .Y(n2814) );
  AND2X4 U2765 ( .A(n2821), .B(n2822), .Y(n2819) );
  OR2X4 U2766 ( .A(n2823), .B(n2824), .Y(n2648) );
  AND2X4 U2767 ( .A(n2825), .B(n2826), .Y(n2824) );
  AND2X4 U2768 ( .A(n2827), .B(n2664), .Y(n2826) );
  OR2X4 U2769 ( .A(n2828), .B(n2829), .Y(n2664) );
  OR2X4 U2770 ( .A(n2830), .B(n2831), .Y(n2827) );
  INVX4 U2771 ( .A(n2663), .Y(n2825) );
  AND2X4 U2772 ( .A(n2663), .B(n2832), .Y(n2823) );
  OR2X4 U2773 ( .A(n2833), .B(n2662), .Y(n2832) );
  AND2X4 U2774 ( .A(n2829), .B(n2828), .Y(n2662) );
  AND2X4 U2775 ( .A(n2830), .B(n2831), .Y(n2833) );
  INVX4 U2776 ( .A(n2828), .Y(n2831) );
  AND2X4 U2777 ( .A(B[1]), .B(A[10]), .Y(n2828) );
  INVX4 U2778 ( .A(n2829), .Y(n2830) );
  OR2X4 U2779 ( .A(n2834), .B(n2835), .Y(n2829) );
  AND2X4 U2780 ( .A(n2836), .B(n2837), .Y(n2834) );
  OR2X4 U2781 ( .A(n2838), .B(n2839), .Y(n2663) );
  AND2X4 U2782 ( .A(n2840), .B(n2841), .Y(n2839) );
  AND2X4 U2783 ( .A(n2842), .B(n2679), .Y(n2841) );
  OR2X4 U2784 ( .A(n2843), .B(n2844), .Y(n2679) );
  OR2X4 U2785 ( .A(n2845), .B(n2846), .Y(n2842) );
  INVX4 U2786 ( .A(n2678), .Y(n2840) );
  AND2X4 U2787 ( .A(n2678), .B(n2847), .Y(n2838) );
  OR2X4 U2788 ( .A(n2848), .B(n2677), .Y(n2847) );
  AND2X4 U2789 ( .A(n2844), .B(n2843), .Y(n2677) );
  AND2X4 U2790 ( .A(n2845), .B(n2846), .Y(n2848) );
  INVX4 U2791 ( .A(n2843), .Y(n2846) );
  AND2X4 U2792 ( .A(B[2]), .B(A[9]), .Y(n2843) );
  INVX4 U2793 ( .A(n2844), .Y(n2845) );
  OR2X4 U2794 ( .A(n2849), .B(n2850), .Y(n2844) );
  AND2X4 U2795 ( .A(n2851), .B(n2852), .Y(n2849) );
  OR2X4 U2796 ( .A(n2853), .B(n2854), .Y(n2678) );
  AND2X4 U2797 ( .A(n2855), .B(n2856), .Y(n2854) );
  AND2X4 U2798 ( .A(n2857), .B(n2694), .Y(n2856) );
  OR2X4 U2799 ( .A(n2858), .B(n2859), .Y(n2694) );
  OR2X4 U2800 ( .A(n2860), .B(n2861), .Y(n2857) );
  INVX4 U2801 ( .A(n2693), .Y(n2855) );
  AND2X4 U2802 ( .A(n2693), .B(n2862), .Y(n2853) );
  OR2X4 U2803 ( .A(n2863), .B(n2692), .Y(n2862) );
  AND2X4 U2804 ( .A(n2859), .B(n2858), .Y(n2692) );
  AND2X4 U2805 ( .A(n2860), .B(n2861), .Y(n2863) );
  INVX4 U2806 ( .A(n2858), .Y(n2861) );
  AND2X4 U2807 ( .A(B[3]), .B(A[8]), .Y(n2858) );
  INVX4 U2808 ( .A(n2859), .Y(n2860) );
  OR2X4 U2809 ( .A(n2864), .B(n2865), .Y(n2859) );
  AND2X4 U2810 ( .A(n2866), .B(n2867), .Y(n2864) );
  OR2X4 U2811 ( .A(n2868), .B(n2869), .Y(n2693) );
  AND2X4 U2812 ( .A(n2870), .B(n2871), .Y(n2869) );
  AND2X4 U2813 ( .A(n2872), .B(n2709), .Y(n2871) );
  OR2X4 U2814 ( .A(n2873), .B(n2874), .Y(n2709) );
  OR2X4 U2815 ( .A(n2875), .B(n2876), .Y(n2872) );
  INVX4 U2816 ( .A(n2708), .Y(n2870) );
  AND2X4 U2817 ( .A(n2708), .B(n2877), .Y(n2868) );
  OR2X4 U2818 ( .A(n2878), .B(n2707), .Y(n2877) );
  AND2X4 U2819 ( .A(n2874), .B(n2873), .Y(n2707) );
  AND2X4 U2820 ( .A(n2875), .B(n2876), .Y(n2878) );
  INVX4 U2821 ( .A(n2873), .Y(n2876) );
  AND2X4 U2822 ( .A(B[4]), .B(A[7]), .Y(n2873) );
  INVX4 U2823 ( .A(n2874), .Y(n2875) );
  OR2X4 U2824 ( .A(n2879), .B(n2880), .Y(n2874) );
  AND2X4 U2825 ( .A(n2881), .B(n2882), .Y(n2879) );
  OR2X4 U2826 ( .A(n2883), .B(n2884), .Y(n2708) );
  AND2X4 U2827 ( .A(n2885), .B(n2886), .Y(n2884) );
  AND2X4 U2828 ( .A(n2887), .B(n2724), .Y(n2886) );
  OR2X4 U2829 ( .A(n2888), .B(n2889), .Y(n2724) );
  OR2X4 U2830 ( .A(n2890), .B(n2891), .Y(n2887) );
  INVX4 U2831 ( .A(n2723), .Y(n2885) );
  AND2X4 U2832 ( .A(n2723), .B(n2892), .Y(n2883) );
  OR2X4 U2833 ( .A(n2893), .B(n2722), .Y(n2892) );
  AND2X4 U2834 ( .A(n2889), .B(n2888), .Y(n2722) );
  AND2X4 U2835 ( .A(n2890), .B(n2891), .Y(n2893) );
  INVX4 U2836 ( .A(n2888), .Y(n2891) );
  AND2X4 U2837 ( .A(B[5]), .B(A[6]), .Y(n2888) );
  INVX4 U2838 ( .A(n2889), .Y(n2890) );
  OR2X4 U2839 ( .A(n2894), .B(n2895), .Y(n2889) );
  AND2X4 U2840 ( .A(n2896), .B(n2897), .Y(n2894) );
  OR2X4 U2841 ( .A(n2898), .B(n2899), .Y(n2723) );
  AND2X4 U2842 ( .A(n2900), .B(n2901), .Y(n2899) );
  AND2X4 U2843 ( .A(n2902), .B(n2739), .Y(n2901) );
  OR2X4 U2844 ( .A(n2903), .B(n2904), .Y(n2739) );
  OR2X4 U2845 ( .A(n2905), .B(n2906), .Y(n2902) );
  INVX4 U2846 ( .A(n2738), .Y(n2900) );
  AND2X4 U2847 ( .A(n2738), .B(n2907), .Y(n2898) );
  OR2X4 U2848 ( .A(n2908), .B(n2737), .Y(n2907) );
  AND2X4 U2849 ( .A(n2904), .B(n2903), .Y(n2737) );
  AND2X4 U2850 ( .A(n2905), .B(n2906), .Y(n2908) );
  INVX4 U2851 ( .A(n2903), .Y(n2906) );
  AND2X4 U2852 ( .A(B[6]), .B(A[5]), .Y(n2903) );
  INVX4 U2853 ( .A(n2904), .Y(n2905) );
  OR2X4 U2854 ( .A(n2909), .B(n2910), .Y(n2904) );
  AND2X4 U2855 ( .A(n2911), .B(n2912), .Y(n2909) );
  OR2X4 U2856 ( .A(n2913), .B(n2914), .Y(n2738) );
  AND2X4 U2857 ( .A(n2915), .B(n2916), .Y(n2914) );
  AND2X4 U2858 ( .A(n2917), .B(n2754), .Y(n2916) );
  OR2X4 U2859 ( .A(n2918), .B(n2919), .Y(n2754) );
  OR2X4 U2860 ( .A(n2920), .B(n2921), .Y(n2917) );
  INVX4 U2861 ( .A(n2753), .Y(n2915) );
  AND2X4 U2862 ( .A(n2753), .B(n2922), .Y(n2913) );
  OR2X4 U2863 ( .A(n2923), .B(n2752), .Y(n2922) );
  AND2X4 U2864 ( .A(n2919), .B(n2918), .Y(n2752) );
  AND2X4 U2865 ( .A(n2920), .B(n2921), .Y(n2923) );
  INVX4 U2866 ( .A(n2918), .Y(n2921) );
  AND2X4 U2867 ( .A(B[7]), .B(A[4]), .Y(n2918) );
  INVX4 U2868 ( .A(n2919), .Y(n2920) );
  OR2X4 U2869 ( .A(n2924), .B(n2925), .Y(n2919) );
  AND2X4 U2870 ( .A(n2926), .B(n2927), .Y(n2924) );
  OR2X4 U2871 ( .A(n2928), .B(n2929), .Y(n2927) );
  OR2X4 U2872 ( .A(n2930), .B(n2931), .Y(n2753) );
  AND2X4 U2873 ( .A(n2932), .B(n2933), .Y(n2931) );
  INVX4 U2874 ( .A(n2768), .Y(n2933) );
  OR2X4 U2875 ( .A(n2934), .B(n2935), .Y(n2932) );
  AND2X4 U2876 ( .A(n2770), .B(n2936), .Y(n2935) );
  AND2X4 U2877 ( .A(n2771), .B(n2937), .Y(n2934) );
  AND2X4 U2878 ( .A(n2768), .B(n2938), .Y(n2930) );
  OR2X4 U2879 ( .A(n2939), .B(n2767), .Y(n2938) );
  AND2X4 U2880 ( .A(n2770), .B(n2771), .Y(n2767) );
  INVX4 U2881 ( .A(n2936), .Y(n2771) );
  AND2X4 U2882 ( .A(n2937), .B(n2936), .Y(n2939) );
  OR2X4 U2883 ( .A(n2940), .B(n633), .Y(n2936) );
  AND2X4 U2884 ( .A(n2941), .B(n2942), .Y(n2940) );
  OR2X4 U2885 ( .A(n2943), .B(n2783), .Y(n2942) );
  AND2X4 U2886 ( .A(n2024), .B(n2944), .Y(n2943) );
  OR2X4 U2887 ( .A(n2945), .B(n1804), .Y(n2944) );
  OR2X4 U2888 ( .A(n2945), .B(n142), .Y(n2941) );
  INVX4 U2889 ( .A(n2770), .Y(n2937) );
  AND2X4 U2890 ( .A(B[8]), .B(A[3]), .Y(n2770) );
  OR2X4 U2891 ( .A(n2946), .B(n2947), .Y(n2768) );
  AND2X4 U2892 ( .A(n2948), .B(n2788), .Y(n2947) );
  INVX4 U2893 ( .A(n2949), .Y(n2788) );
  AND2X4 U2894 ( .A(B[9]), .B(n2950), .Y(n2948) );
  OR2X4 U2895 ( .A(n131), .B(n2951), .Y(n2950) );
  OR2X4 U2896 ( .A(n2952), .B(n2953), .Y(n2951) );
  AND2X4 U2897 ( .A(n2233), .B(B[10]), .Y(n2953) );
  AND2X4 U2898 ( .A(A[2]), .B(n423), .Y(n2952) );
  AND2X4 U2899 ( .A(n2954), .B(n2949), .Y(n2946) );
  OR2X4 U2900 ( .A(n2955), .B(n2956), .Y(n2949) );
  AND2X4 U2901 ( .A(B[11]), .B(n2957), .Y(n2956) );
  OR2X4 U2902 ( .A(n2958), .B(n1207), .Y(n2957) );
  AND2X4 U2903 ( .A(A[0]), .B(n423), .Y(n2958) );
  AND2X4 U2904 ( .A(B[10]), .B(n2959), .Y(n2955) );
  OR2X4 U2905 ( .A(n2960), .B(n1210), .Y(n2959) );
  AND2X4 U2906 ( .A(A[1]), .B(n2423), .Y(n2960) );
  INVX4 U2907 ( .A(B[11]), .Y(n2423) );
  OR2X4 U2908 ( .A(n2961), .B(n2962), .Y(n2954) );
  OR2X4 U2909 ( .A(n137), .B(n2783), .Y(n2962) );
  OR2X4 U2910 ( .A(n2963), .B(n2964), .Y(n2961) );
  AND2X4 U2911 ( .A(n141), .B(B[10]), .Y(n2964) );
  AND2X4 U2912 ( .A(n142), .B(n423), .Y(n2963) );
  OR2X4 U2913 ( .A(n2965), .B(n2966), .Y(Y[10]) );
  AND2X4 U2914 ( .A(n2967), .B(n2968), .Y(n2966) );
  AND2X4 U2915 ( .A(n2969), .B(n2822), .Y(n2968) );
  OR2X4 U2916 ( .A(n2970), .B(n2971), .Y(n2822) );
  OR2X4 U2917 ( .A(n2972), .B(n2973), .Y(n2969) );
  INVX4 U2918 ( .A(n2821), .Y(n2967) );
  AND2X4 U2919 ( .A(n2821), .B(n2974), .Y(n2965) );
  OR2X4 U2920 ( .A(n2975), .B(n2820), .Y(n2974) );
  AND2X4 U2921 ( .A(n2971), .B(n2970), .Y(n2820) );
  AND2X4 U2922 ( .A(n2972), .B(n2973), .Y(n2975) );
  INVX4 U2923 ( .A(n2970), .Y(n2973) );
  AND2X4 U2924 ( .A(B[0]), .B(A[10]), .Y(n2970) );
  INVX4 U2925 ( .A(n2971), .Y(n2972) );
  OR2X4 U2926 ( .A(n2976), .B(n14), .Y(n2971) );
  AND2X4 U2927 ( .A(n16), .B(n15), .Y(n14) );
  AND2X4 U2928 ( .A(n7), .B(n11), .Y(n2976) );
  OR2X4 U2929 ( .A(n2977), .B(n2978), .Y(n11) );
  OR2X4 U2930 ( .A(n2979), .B(n2980), .Y(n2978) );
  AND2X4 U2931 ( .A(n2981), .B(n2982), .Y(n2980) );
  INVX4 U2932 ( .A(n2983), .Y(n2982) );
  AND2X4 U2933 ( .A(n2984), .B(n2985), .Y(n2981) );
  OR2X4 U2934 ( .A(n2986), .B(n2987), .Y(n2985) );
  OR2X4 U2935 ( .A(n2988), .B(n2989), .Y(n2984) );
  AND2X4 U2936 ( .A(n2990), .B(n2983), .Y(n2979) );
  AND2X4 U2937 ( .A(n2988), .B(n2989), .Y(n2990) );
  INVX4 U2938 ( .A(n2986), .Y(n2989) );
  INVX4 U2939 ( .A(n2987), .Y(n2988) );
  AND2X4 U2940 ( .A(n2991), .B(n2987), .Y(n2977) );
  OR2X4 U2941 ( .A(n15), .B(n16), .Y(n7) );
  OR2X4 U2942 ( .A(n2992), .B(n28), .Y(n16) );
  AND2X4 U2943 ( .A(n30), .B(n29), .Y(n28) );
  AND2X4 U2944 ( .A(n22), .B(n25), .Y(n2992) );
  OR2X4 U2945 ( .A(n2993), .B(n2994), .Y(n25) );
  OR2X4 U2946 ( .A(n2995), .B(n2996), .Y(n2994) );
  AND2X4 U2947 ( .A(n2997), .B(n2998), .Y(n2996) );
  INVX4 U2948 ( .A(n2999), .Y(n2998) );
  AND2X4 U2949 ( .A(n3000), .B(n3001), .Y(n2997) );
  OR2X4 U2950 ( .A(n3002), .B(n3003), .Y(n3001) );
  OR2X4 U2951 ( .A(n3004), .B(n3005), .Y(n3000) );
  AND2X4 U2952 ( .A(n3006), .B(n2999), .Y(n2995) );
  AND2X4 U2953 ( .A(n3004), .B(n3005), .Y(n3006) );
  INVX4 U2954 ( .A(n3002), .Y(n3005) );
  INVX4 U2955 ( .A(n3003), .Y(n3004) );
  AND2X4 U2956 ( .A(n3007), .B(n3003), .Y(n2993) );
  OR2X4 U2957 ( .A(n29), .B(n30), .Y(n22) );
  OR2X4 U2958 ( .A(n3008), .B(n42), .Y(n30) );
  AND2X4 U2959 ( .A(n44), .B(n43), .Y(n42) );
  AND2X4 U2960 ( .A(n36), .B(n39), .Y(n3008) );
  OR2X4 U2961 ( .A(n3009), .B(n3010), .Y(n39) );
  OR2X4 U2962 ( .A(n3011), .B(n3012), .Y(n3010) );
  AND2X4 U2963 ( .A(n3013), .B(n3014), .Y(n3012) );
  INVX4 U2964 ( .A(n3015), .Y(n3014) );
  AND2X4 U2965 ( .A(n3016), .B(n3017), .Y(n3013) );
  OR2X4 U2966 ( .A(n3018), .B(n3019), .Y(n3017) );
  OR2X4 U2967 ( .A(n3020), .B(n3021), .Y(n3016) );
  AND2X4 U2968 ( .A(n3022), .B(n3015), .Y(n3011) );
  AND2X4 U2969 ( .A(n3020), .B(n3021), .Y(n3022) );
  INVX4 U2970 ( .A(n3018), .Y(n3021) );
  INVX4 U2971 ( .A(n3019), .Y(n3020) );
  AND2X4 U2972 ( .A(n3023), .B(n3019), .Y(n3009) );
  OR2X4 U2973 ( .A(n43), .B(n44), .Y(n36) );
  OR2X4 U2974 ( .A(n3024), .B(n56), .Y(n44) );
  AND2X4 U2975 ( .A(n58), .B(n57), .Y(n56) );
  AND2X4 U2976 ( .A(n50), .B(n53), .Y(n3024) );
  OR2X4 U2977 ( .A(n3025), .B(n3026), .Y(n53) );
  OR2X4 U2978 ( .A(n3027), .B(n3028), .Y(n3026) );
  AND2X4 U2979 ( .A(n3029), .B(n3030), .Y(n3028) );
  INVX4 U2980 ( .A(n3031), .Y(n3030) );
  AND2X4 U2981 ( .A(n3032), .B(n3033), .Y(n3029) );
  OR2X4 U2982 ( .A(n3034), .B(n3035), .Y(n3033) );
  OR2X4 U2983 ( .A(n3036), .B(n3037), .Y(n3032) );
  AND2X4 U2984 ( .A(n3038), .B(n3031), .Y(n3027) );
  AND2X4 U2985 ( .A(n3036), .B(n3037), .Y(n3038) );
  INVX4 U2986 ( .A(n3034), .Y(n3037) );
  INVX4 U2987 ( .A(n3035), .Y(n3036) );
  AND2X4 U2988 ( .A(n3039), .B(n3035), .Y(n3025) );
  OR2X4 U2989 ( .A(n57), .B(n58), .Y(n50) );
  OR2X4 U2990 ( .A(n3040), .B(n70), .Y(n58) );
  AND2X4 U2991 ( .A(n72), .B(n71), .Y(n70) );
  AND2X4 U2992 ( .A(n64), .B(n67), .Y(n3040) );
  OR2X4 U2993 ( .A(n3041), .B(n3042), .Y(n67) );
  OR2X4 U2994 ( .A(n3043), .B(n3044), .Y(n3042) );
  AND2X4 U2995 ( .A(n3045), .B(n3046), .Y(n3044) );
  INVX4 U2996 ( .A(n3047), .Y(n3046) );
  AND2X4 U2997 ( .A(n3048), .B(n3049), .Y(n3045) );
  OR2X4 U2998 ( .A(n3050), .B(n3051), .Y(n3049) );
  OR2X4 U2999 ( .A(n3052), .B(n3053), .Y(n3048) );
  AND2X4 U3000 ( .A(n3054), .B(n3047), .Y(n3043) );
  AND2X4 U3001 ( .A(n3052), .B(n3053), .Y(n3054) );
  INVX4 U3002 ( .A(n3050), .Y(n3053) );
  INVX4 U3003 ( .A(n3051), .Y(n3052) );
  AND2X4 U3004 ( .A(n3055), .B(n3051), .Y(n3041) );
  OR2X4 U3005 ( .A(n71), .B(n72), .Y(n64) );
  OR2X4 U3006 ( .A(n3056), .B(n84), .Y(n72) );
  AND2X4 U3007 ( .A(n86), .B(n85), .Y(n84) );
  AND2X4 U3008 ( .A(n78), .B(n81), .Y(n3056) );
  OR2X4 U3009 ( .A(n3057), .B(n3058), .Y(n81) );
  OR2X4 U3010 ( .A(n3059), .B(n3060), .Y(n3058) );
  AND2X4 U3011 ( .A(n3061), .B(n3062), .Y(n3060) );
  INVX4 U3012 ( .A(n3063), .Y(n3062) );
  OR2X4 U3013 ( .A(n3064), .B(n3065), .Y(n3061) );
  AND2X4 U3014 ( .A(n3066), .B(n3067), .Y(n3065) );
  AND2X4 U3015 ( .A(n3068), .B(n3069), .Y(n3064) );
  AND2X4 U3016 ( .A(n3070), .B(n3063), .Y(n3059) );
  AND2X4 U3017 ( .A(n3069), .B(n3067), .Y(n3070) );
  INVX4 U3018 ( .A(n3066), .Y(n3069) );
  AND2X4 U3019 ( .A(n3071), .B(n3068), .Y(n3057) );
  OR2X4 U3020 ( .A(n85), .B(n86), .Y(n78) );
  OR2X4 U3021 ( .A(n3072), .B(n98), .Y(n86) );
  AND2X4 U3022 ( .A(n100), .B(n99), .Y(n98) );
  AND2X4 U3023 ( .A(n95), .B(n92), .Y(n3072) );
  OR2X4 U3024 ( .A(n99), .B(n100), .Y(n92) );
  OR2X4 U3025 ( .A(n3073), .B(n3074), .Y(n100) );
  AND2X4 U3026 ( .A(n3075), .B(B[0]), .Y(n3074) );
  AND2X4 U3027 ( .A(A[2]), .B(n134), .Y(n3075) );
  AND2X4 U3028 ( .A(n3076), .B(Y[0]), .Y(n3073) );
  AND2X4 U3029 ( .A(n145), .B(n3077), .Y(n3076) );
  INVX4 U3030 ( .A(n144), .Y(n3077) );
  AND2X4 U3031 ( .A(n142), .B(n128), .Y(n144) );
  INVX4 U3032 ( .A(n134), .Y(n128) );
  OR2X4 U3033 ( .A(n3078), .B(n3079), .Y(n134) );
  OR2X4 U3034 ( .A(n3080), .B(n3081), .Y(n3079) );
  AND2X4 U3035 ( .A(B[2]), .B(n3082), .Y(n3081) );
  OR2X4 U3036 ( .A(n3083), .B(n1207), .Y(n3082) );
  AND2X4 U3037 ( .A(A[0]), .B(n132), .Y(n3083) );
  AND2X4 U3038 ( .A(n145), .B(n1622), .Y(n3080) );
  AND2X4 U3039 ( .A(n1210), .B(B[1]), .Y(n3078) );
  AND2X4 U3040 ( .A(A[1]), .B(B[1]), .Y(n145) );
  AND2X4 U3041 ( .A(A[3]), .B(B[0]), .Y(n99) );
  OR2X4 U3042 ( .A(n3084), .B(n3085), .Y(n95) );
  AND2X4 U3043 ( .A(n3086), .B(n3087), .Y(n3085) );
  AND2X4 U3044 ( .A(B[1]), .B(n3088), .Y(n3086) );
  OR2X4 U3045 ( .A(n131), .B(n3089), .Y(n3088) );
  OR2X4 U3046 ( .A(n3090), .B(n3091), .Y(n3089) );
  AND2X4 U3047 ( .A(n2233), .B(B[2]), .Y(n3091) );
  AND2X4 U3048 ( .A(A[2]), .B(n1622), .Y(n3090) );
  AND2X4 U3049 ( .A(n3092), .B(n3093), .Y(n3084) );
  OR2X4 U3050 ( .A(n3094), .B(n3095), .Y(n3092) );
  OR2X4 U3051 ( .A(n137), .B(n132), .Y(n3095) );
  OR2X4 U3052 ( .A(n3096), .B(n3097), .Y(n3094) );
  AND2X4 U3053 ( .A(n141), .B(B[2]), .Y(n3097) );
  AND2X4 U3054 ( .A(n142), .B(n1622), .Y(n3096) );
  AND2X4 U3055 ( .A(A[4]), .B(B[0]), .Y(n85) );
  AND2X4 U3056 ( .A(A[5]), .B(B[0]), .Y(n71) );
  AND2X4 U3057 ( .A(A[6]), .B(B[0]), .Y(n57) );
  AND2X4 U3058 ( .A(A[7]), .B(B[0]), .Y(n43) );
  AND2X4 U3059 ( .A(A[8]), .B(B[0]), .Y(n29) );
  AND2X4 U3060 ( .A(A[9]), .B(B[0]), .Y(n15) );
  OR2X4 U3061 ( .A(n3098), .B(n3099), .Y(n2821) );
  AND2X4 U3062 ( .A(n3100), .B(n3101), .Y(n3099) );
  AND2X4 U3063 ( .A(n3102), .B(n2837), .Y(n3101) );
  OR2X4 U3064 ( .A(n3103), .B(n3104), .Y(n2837) );
  OR2X4 U3065 ( .A(n3105), .B(n3106), .Y(n3102) );
  INVX4 U3066 ( .A(n2836), .Y(n3100) );
  AND2X4 U3067 ( .A(n2836), .B(n3107), .Y(n3098) );
  OR2X4 U3068 ( .A(n3108), .B(n2835), .Y(n3107) );
  AND2X4 U3069 ( .A(n3104), .B(n3103), .Y(n2835) );
  AND2X4 U3070 ( .A(n3105), .B(n3106), .Y(n3108) );
  INVX4 U3071 ( .A(n3103), .Y(n3106) );
  AND2X4 U3072 ( .A(B[1]), .B(A[9]), .Y(n3103) );
  INVX4 U3073 ( .A(n3104), .Y(n3105) );
  OR2X4 U3074 ( .A(n3109), .B(n2991), .Y(n3104) );
  AND2X4 U3075 ( .A(n2983), .B(n2986), .Y(n2991) );
  AND2X4 U3076 ( .A(n3110), .B(n2987), .Y(n3109) );
  OR2X4 U3077 ( .A(n3111), .B(n3007), .Y(n2987) );
  AND2X4 U3078 ( .A(n2999), .B(n3002), .Y(n3007) );
  AND2X4 U3079 ( .A(n3112), .B(n3003), .Y(n3111) );
  OR2X4 U3080 ( .A(n3113), .B(n3023), .Y(n3003) );
  AND2X4 U3081 ( .A(n3015), .B(n3018), .Y(n3023) );
  AND2X4 U3082 ( .A(n3114), .B(n3019), .Y(n3113) );
  OR2X4 U3083 ( .A(n3115), .B(n3039), .Y(n3019) );
  AND2X4 U3084 ( .A(n3031), .B(n3034), .Y(n3039) );
  AND2X4 U3085 ( .A(n3116), .B(n3035), .Y(n3115) );
  OR2X4 U3086 ( .A(n3117), .B(n3055), .Y(n3035) );
  AND2X4 U3087 ( .A(n3047), .B(n3050), .Y(n3055) );
  AND2X4 U3088 ( .A(n3118), .B(n3051), .Y(n3117) );
  OR2X4 U3089 ( .A(n3119), .B(n3071), .Y(n3051) );
  AND2X4 U3090 ( .A(n3063), .B(n3066), .Y(n3071) );
  AND2X4 U3091 ( .A(n3068), .B(n3120), .Y(n3119) );
  OR2X4 U3092 ( .A(n3066), .B(n3063), .Y(n3120) );
  OR2X4 U3093 ( .A(n3121), .B(n3122), .Y(n3063) );
  AND2X4 U3094 ( .A(n3123), .B(n3124), .Y(n3122) );
  AND2X4 U3095 ( .A(B[2]), .B(n3125), .Y(n3123) );
  OR2X4 U3096 ( .A(n131), .B(n3126), .Y(n3125) );
  OR2X4 U3097 ( .A(n3127), .B(n3128), .Y(n3126) );
  AND2X4 U3098 ( .A(n2233), .B(B[3]), .Y(n3128) );
  AND2X4 U3099 ( .A(A[2]), .B(n3129), .Y(n3127) );
  AND2X4 U3100 ( .A(n3130), .B(n3131), .Y(n3121) );
  OR2X4 U3101 ( .A(n3132), .B(n3133), .Y(n3130) );
  OR2X4 U3102 ( .A(n137), .B(n1622), .Y(n3133) );
  OR2X4 U3103 ( .A(n3134), .B(n3135), .Y(n3132) );
  AND2X4 U3104 ( .A(n141), .B(B[3]), .Y(n3135) );
  AND2X4 U3105 ( .A(n142), .B(n3129), .Y(n3134) );
  AND2X4 U3106 ( .A(A[3]), .B(B[1]), .Y(n3066) );
  INVX4 U3107 ( .A(n3067), .Y(n3068) );
  OR2X4 U3108 ( .A(n3136), .B(n132), .Y(n3067) );
  INVX4 U3109 ( .A(B[1]), .Y(n132) );
  AND2X4 U3110 ( .A(n3137), .B(n3138), .Y(n3136) );
  OR2X4 U3111 ( .A(n3139), .B(n1622), .Y(n3138) );
  AND2X4 U3112 ( .A(n2024), .B(n3140), .Y(n3139) );
  OR2X4 U3113 ( .A(n3087), .B(n1804), .Y(n3140) );
  OR2X4 U3114 ( .A(n3087), .B(n142), .Y(n3137) );
  INVX4 U3115 ( .A(n3093), .Y(n3087) );
  OR2X4 U3116 ( .A(n3141), .B(n3142), .Y(n3093) );
  AND2X4 U3117 ( .A(B[3]), .B(n3143), .Y(n3142) );
  OR2X4 U3118 ( .A(n3144), .B(n1207), .Y(n3143) );
  AND2X4 U3119 ( .A(A[0]), .B(n1622), .Y(n3144) );
  AND2X4 U3120 ( .A(B[2]), .B(n3145), .Y(n3141) );
  OR2X4 U3121 ( .A(n3146), .B(n1210), .Y(n3145) );
  AND2X4 U3122 ( .A(A[1]), .B(n3129), .Y(n3146) );
  OR2X4 U3123 ( .A(n3050), .B(n3047), .Y(n3118) );
  OR2X4 U3124 ( .A(n3147), .B(n3148), .Y(n3047) );
  OR2X4 U3125 ( .A(n3149), .B(n3150), .Y(n3148) );
  AND2X4 U3126 ( .A(n3151), .B(n3152), .Y(n3150) );
  INVX4 U3127 ( .A(n3153), .Y(n3152) );
  OR2X4 U3128 ( .A(n3154), .B(n3155), .Y(n3151) );
  AND2X4 U3129 ( .A(n3156), .B(n3157), .Y(n3155) );
  AND2X4 U3130 ( .A(n3158), .B(n3159), .Y(n3154) );
  AND2X4 U3131 ( .A(n3160), .B(n3153), .Y(n3149) );
  AND2X4 U3132 ( .A(n3159), .B(n3157), .Y(n3160) );
  INVX4 U3133 ( .A(n3156), .Y(n3159) );
  AND2X4 U3134 ( .A(n3161), .B(n3158), .Y(n3147) );
  AND2X4 U3135 ( .A(A[4]), .B(B[1]), .Y(n3050) );
  OR2X4 U3136 ( .A(n3034), .B(n3031), .Y(n3116) );
  OR2X4 U3137 ( .A(n3162), .B(n3163), .Y(n3031) );
  OR2X4 U3138 ( .A(n3164), .B(n3165), .Y(n3163) );
  AND2X4 U3139 ( .A(n3166), .B(n3167), .Y(n3165) );
  INVX4 U3140 ( .A(n3168), .Y(n3167) );
  AND2X4 U3141 ( .A(n3169), .B(n3170), .Y(n3166) );
  OR2X4 U3142 ( .A(n3171), .B(n3172), .Y(n3170) );
  OR2X4 U3143 ( .A(n3173), .B(n3174), .Y(n3169) );
  AND2X4 U3144 ( .A(n3175), .B(n3168), .Y(n3164) );
  AND2X4 U3145 ( .A(n3173), .B(n3174), .Y(n3175) );
  INVX4 U3146 ( .A(n3171), .Y(n3174) );
  INVX4 U3147 ( .A(n3172), .Y(n3173) );
  AND2X4 U3148 ( .A(n3176), .B(n3172), .Y(n3162) );
  AND2X4 U3149 ( .A(A[5]), .B(B[1]), .Y(n3034) );
  OR2X4 U3150 ( .A(n3018), .B(n3015), .Y(n3114) );
  OR2X4 U3151 ( .A(n3177), .B(n3178), .Y(n3015) );
  OR2X4 U3152 ( .A(n3179), .B(n3180), .Y(n3178) );
  AND2X4 U3153 ( .A(n3181), .B(n3182), .Y(n3180) );
  INVX4 U3154 ( .A(n3183), .Y(n3182) );
  AND2X4 U3155 ( .A(n3184), .B(n3185), .Y(n3181) );
  OR2X4 U3156 ( .A(n3186), .B(n3187), .Y(n3185) );
  OR2X4 U3157 ( .A(n3188), .B(n3189), .Y(n3184) );
  AND2X4 U3158 ( .A(n3190), .B(n3183), .Y(n3179) );
  AND2X4 U3159 ( .A(n3188), .B(n3189), .Y(n3190) );
  INVX4 U3160 ( .A(n3186), .Y(n3189) );
  INVX4 U3161 ( .A(n3187), .Y(n3188) );
  AND2X4 U3162 ( .A(n3191), .B(n3187), .Y(n3177) );
  AND2X4 U3163 ( .A(A[6]), .B(B[1]), .Y(n3018) );
  OR2X4 U3164 ( .A(n3002), .B(n2999), .Y(n3112) );
  OR2X4 U3165 ( .A(n3192), .B(n3193), .Y(n2999) );
  OR2X4 U3166 ( .A(n3194), .B(n3195), .Y(n3193) );
  AND2X4 U3167 ( .A(n3196), .B(n3197), .Y(n3195) );
  INVX4 U3168 ( .A(n3198), .Y(n3197) );
  AND2X4 U3169 ( .A(n3199), .B(n3200), .Y(n3196) );
  OR2X4 U3170 ( .A(n3201), .B(n3202), .Y(n3200) );
  OR2X4 U3171 ( .A(n3203), .B(n3204), .Y(n3199) );
  AND2X4 U3172 ( .A(n3205), .B(n3198), .Y(n3194) );
  AND2X4 U3173 ( .A(n3203), .B(n3204), .Y(n3205) );
  INVX4 U3174 ( .A(n3201), .Y(n3204) );
  INVX4 U3175 ( .A(n3202), .Y(n3203) );
  AND2X4 U3176 ( .A(n3206), .B(n3202), .Y(n3192) );
  AND2X4 U3177 ( .A(A[7]), .B(B[1]), .Y(n3002) );
  OR2X4 U3178 ( .A(n2986), .B(n2983), .Y(n3110) );
  OR2X4 U3179 ( .A(n3207), .B(n3208), .Y(n2983) );
  OR2X4 U3180 ( .A(n3209), .B(n3210), .Y(n3208) );
  AND2X4 U3181 ( .A(n3211), .B(n3212), .Y(n3210) );
  INVX4 U3182 ( .A(n3213), .Y(n3212) );
  AND2X4 U3183 ( .A(n3214), .B(n3215), .Y(n3211) );
  OR2X4 U3184 ( .A(n3216), .B(n3217), .Y(n3215) );
  OR2X4 U3185 ( .A(n3218), .B(n3219), .Y(n3214) );
  AND2X4 U3186 ( .A(n3220), .B(n3213), .Y(n3209) );
  AND2X4 U3187 ( .A(n3218), .B(n3219), .Y(n3220) );
  INVX4 U3188 ( .A(n3216), .Y(n3219) );
  INVX4 U3189 ( .A(n3217), .Y(n3218) );
  AND2X4 U3190 ( .A(n3221), .B(n3217), .Y(n3207) );
  AND2X4 U3191 ( .A(B[1]), .B(A[8]), .Y(n2986) );
  OR2X4 U3192 ( .A(n3222), .B(n3223), .Y(n2836) );
  AND2X4 U3193 ( .A(n3224), .B(n3225), .Y(n3223) );
  AND2X4 U3194 ( .A(n3226), .B(n2852), .Y(n3225) );
  OR2X4 U3195 ( .A(n3227), .B(n3228), .Y(n2852) );
  OR2X4 U3196 ( .A(n3229), .B(n3230), .Y(n3226) );
  INVX4 U3197 ( .A(n2851), .Y(n3224) );
  AND2X4 U3198 ( .A(n2851), .B(n3231), .Y(n3222) );
  OR2X4 U3199 ( .A(n3232), .B(n2850), .Y(n3231) );
  AND2X4 U3200 ( .A(n3228), .B(n3227), .Y(n2850) );
  AND2X4 U3201 ( .A(n3229), .B(n3230), .Y(n3232) );
  INVX4 U3202 ( .A(n3227), .Y(n3230) );
  AND2X4 U3203 ( .A(B[2]), .B(A[8]), .Y(n3227) );
  INVX4 U3204 ( .A(n3228), .Y(n3229) );
  OR2X4 U3205 ( .A(n3233), .B(n3221), .Y(n3228) );
  AND2X4 U3206 ( .A(n3213), .B(n3216), .Y(n3221) );
  AND2X4 U3207 ( .A(n3234), .B(n3217), .Y(n3233) );
  OR2X4 U3208 ( .A(n3235), .B(n3206), .Y(n3217) );
  AND2X4 U3209 ( .A(n3198), .B(n3201), .Y(n3206) );
  AND2X4 U3210 ( .A(n3236), .B(n3202), .Y(n3235) );
  OR2X4 U3211 ( .A(n3237), .B(n3191), .Y(n3202) );
  AND2X4 U3212 ( .A(n3183), .B(n3186), .Y(n3191) );
  AND2X4 U3213 ( .A(n3238), .B(n3187), .Y(n3237) );
  OR2X4 U3214 ( .A(n3239), .B(n3176), .Y(n3187) );
  AND2X4 U3215 ( .A(n3168), .B(n3171), .Y(n3176) );
  AND2X4 U3216 ( .A(n3240), .B(n3172), .Y(n3239) );
  OR2X4 U3217 ( .A(n3241), .B(n3161), .Y(n3172) );
  AND2X4 U3218 ( .A(n3153), .B(n3156), .Y(n3161) );
  AND2X4 U3219 ( .A(n3158), .B(n3242), .Y(n3241) );
  OR2X4 U3220 ( .A(n3156), .B(n3153), .Y(n3242) );
  OR2X4 U3221 ( .A(n3243), .B(n3244), .Y(n3153) );
  AND2X4 U3222 ( .A(n3245), .B(n3246), .Y(n3244) );
  AND2X4 U3223 ( .A(B[3]), .B(n3247), .Y(n3245) );
  OR2X4 U3224 ( .A(n131), .B(n3248), .Y(n3247) );
  OR2X4 U3225 ( .A(n3249), .B(n3250), .Y(n3248) );
  AND2X4 U3226 ( .A(n2233), .B(B[4]), .Y(n3250) );
  AND2X4 U3227 ( .A(A[2]), .B(n1241), .Y(n3249) );
  AND2X4 U3228 ( .A(n3251), .B(n3252), .Y(n3243) );
  OR2X4 U3229 ( .A(n3253), .B(n3254), .Y(n3251) );
  OR2X4 U3230 ( .A(n137), .B(n3129), .Y(n3254) );
  OR2X4 U3231 ( .A(n3255), .B(n3256), .Y(n3253) );
  AND2X4 U3232 ( .A(n141), .B(B[4]), .Y(n3256) );
  AND2X4 U3233 ( .A(n142), .B(n1241), .Y(n3255) );
  AND2X4 U3234 ( .A(A[3]), .B(B[2]), .Y(n3156) );
  INVX4 U3235 ( .A(n3157), .Y(n3158) );
  OR2X4 U3236 ( .A(n3257), .B(n1622), .Y(n3157) );
  INVX4 U3237 ( .A(B[2]), .Y(n1622) );
  AND2X4 U3238 ( .A(n3258), .B(n3259), .Y(n3257) );
  OR2X4 U3239 ( .A(n3260), .B(n3129), .Y(n3259) );
  AND2X4 U3240 ( .A(n2024), .B(n3261), .Y(n3260) );
  OR2X4 U3241 ( .A(n3124), .B(n1804), .Y(n3261) );
  OR2X4 U3242 ( .A(n3124), .B(n142), .Y(n3258) );
  INVX4 U3243 ( .A(n3131), .Y(n3124) );
  OR2X4 U3244 ( .A(n3262), .B(n3263), .Y(n3131) );
  AND2X4 U3245 ( .A(B[4]), .B(n3264), .Y(n3263) );
  OR2X4 U3246 ( .A(n3265), .B(n1207), .Y(n3264) );
  AND2X4 U3247 ( .A(A[0]), .B(n3129), .Y(n3265) );
  AND2X4 U3248 ( .A(B[3]), .B(n3266), .Y(n3262) );
  OR2X4 U3249 ( .A(n3267), .B(n1210), .Y(n3266) );
  AND2X4 U3250 ( .A(A[1]), .B(n1241), .Y(n3267) );
  OR2X4 U3251 ( .A(n3171), .B(n3168), .Y(n3240) );
  OR2X4 U3252 ( .A(n3268), .B(n3269), .Y(n3168) );
  OR2X4 U3253 ( .A(n3270), .B(n3271), .Y(n3269) );
  AND2X4 U3254 ( .A(n3272), .B(n3273), .Y(n3271) );
  INVX4 U3255 ( .A(n3274), .Y(n3273) );
  OR2X4 U3256 ( .A(n3275), .B(n3276), .Y(n3272) );
  AND2X4 U3257 ( .A(n3277), .B(n3278), .Y(n3276) );
  AND2X4 U3258 ( .A(n3279), .B(n3280), .Y(n3275) );
  AND2X4 U3259 ( .A(n3281), .B(n3274), .Y(n3270) );
  AND2X4 U3260 ( .A(n3280), .B(n3278), .Y(n3281) );
  INVX4 U3261 ( .A(n3277), .Y(n3280) );
  AND2X4 U3262 ( .A(n3282), .B(n3279), .Y(n3268) );
  AND2X4 U3263 ( .A(A[4]), .B(B[2]), .Y(n3171) );
  OR2X4 U3264 ( .A(n3186), .B(n3183), .Y(n3238) );
  OR2X4 U3265 ( .A(n3283), .B(n3284), .Y(n3183) );
  OR2X4 U3266 ( .A(n3285), .B(n3286), .Y(n3284) );
  AND2X4 U3267 ( .A(n3287), .B(n3288), .Y(n3286) );
  INVX4 U3268 ( .A(n3289), .Y(n3288) );
  AND2X4 U3269 ( .A(n3290), .B(n3291), .Y(n3287) );
  OR2X4 U3270 ( .A(n3292), .B(n3293), .Y(n3291) );
  OR2X4 U3271 ( .A(n3294), .B(n3295), .Y(n3290) );
  AND2X4 U3272 ( .A(n3296), .B(n3289), .Y(n3285) );
  AND2X4 U3273 ( .A(n3294), .B(n3295), .Y(n3296) );
  INVX4 U3274 ( .A(n3292), .Y(n3295) );
  INVX4 U3275 ( .A(n3293), .Y(n3294) );
  AND2X4 U3276 ( .A(n3297), .B(n3293), .Y(n3283) );
  AND2X4 U3277 ( .A(A[5]), .B(B[2]), .Y(n3186) );
  OR2X4 U3278 ( .A(n3201), .B(n3198), .Y(n3236) );
  OR2X4 U3279 ( .A(n3298), .B(n3299), .Y(n3198) );
  OR2X4 U3280 ( .A(n3300), .B(n3301), .Y(n3299) );
  AND2X4 U3281 ( .A(n3302), .B(n3303), .Y(n3301) );
  INVX4 U3282 ( .A(n3304), .Y(n3303) );
  AND2X4 U3283 ( .A(n3305), .B(n3306), .Y(n3302) );
  OR2X4 U3284 ( .A(n3307), .B(n3308), .Y(n3306) );
  OR2X4 U3285 ( .A(n3309), .B(n3310), .Y(n3305) );
  AND2X4 U3286 ( .A(n3311), .B(n3304), .Y(n3300) );
  AND2X4 U3287 ( .A(n3309), .B(n3310), .Y(n3311) );
  INVX4 U3288 ( .A(n3307), .Y(n3310) );
  INVX4 U3289 ( .A(n3308), .Y(n3309) );
  AND2X4 U3290 ( .A(n3312), .B(n3308), .Y(n3298) );
  AND2X4 U3291 ( .A(A[6]), .B(B[2]), .Y(n3201) );
  OR2X4 U3292 ( .A(n3216), .B(n3213), .Y(n3234) );
  OR2X4 U3293 ( .A(n3313), .B(n3314), .Y(n3213) );
  OR2X4 U3294 ( .A(n3315), .B(n3316), .Y(n3314) );
  AND2X4 U3295 ( .A(n3317), .B(n3318), .Y(n3316) );
  INVX4 U3296 ( .A(n3319), .Y(n3318) );
  AND2X4 U3297 ( .A(n3320), .B(n3321), .Y(n3317) );
  OR2X4 U3298 ( .A(n3322), .B(n3323), .Y(n3321) );
  OR2X4 U3299 ( .A(n3324), .B(n3325), .Y(n3320) );
  AND2X4 U3300 ( .A(n3326), .B(n3319), .Y(n3315) );
  AND2X4 U3301 ( .A(n3324), .B(n3325), .Y(n3326) );
  INVX4 U3302 ( .A(n3322), .Y(n3325) );
  INVX4 U3303 ( .A(n3323), .Y(n3324) );
  AND2X4 U3304 ( .A(n3327), .B(n3323), .Y(n3313) );
  AND2X4 U3305 ( .A(B[2]), .B(A[7]), .Y(n3216) );
  OR2X4 U3306 ( .A(n3328), .B(n3329), .Y(n2851) );
  AND2X4 U3307 ( .A(n3330), .B(n3331), .Y(n3329) );
  AND2X4 U3308 ( .A(n3332), .B(n2867), .Y(n3331) );
  OR2X4 U3309 ( .A(n3333), .B(n3334), .Y(n2867) );
  OR2X4 U3310 ( .A(n3335), .B(n3336), .Y(n3332) );
  INVX4 U3311 ( .A(n2866), .Y(n3330) );
  AND2X4 U3312 ( .A(n2866), .B(n3337), .Y(n3328) );
  OR2X4 U3313 ( .A(n3338), .B(n2865), .Y(n3337) );
  AND2X4 U3314 ( .A(n3334), .B(n3333), .Y(n2865) );
  AND2X4 U3315 ( .A(n3335), .B(n3336), .Y(n3338) );
  INVX4 U3316 ( .A(n3333), .Y(n3336) );
  AND2X4 U3317 ( .A(B[3]), .B(A[7]), .Y(n3333) );
  INVX4 U3318 ( .A(n3334), .Y(n3335) );
  OR2X4 U3319 ( .A(n3339), .B(n3327), .Y(n3334) );
  AND2X4 U3320 ( .A(n3319), .B(n3322), .Y(n3327) );
  AND2X4 U3321 ( .A(n3340), .B(n3323), .Y(n3339) );
  OR2X4 U3322 ( .A(n3341), .B(n3312), .Y(n3323) );
  AND2X4 U3323 ( .A(n3304), .B(n3307), .Y(n3312) );
  AND2X4 U3324 ( .A(n3342), .B(n3308), .Y(n3341) );
  OR2X4 U3325 ( .A(n3343), .B(n3297), .Y(n3308) );
  AND2X4 U3326 ( .A(n3289), .B(n3292), .Y(n3297) );
  AND2X4 U3327 ( .A(n3344), .B(n3293), .Y(n3343) );
  OR2X4 U3328 ( .A(n3345), .B(n3282), .Y(n3293) );
  AND2X4 U3329 ( .A(n3274), .B(n3277), .Y(n3282) );
  AND2X4 U3330 ( .A(n3279), .B(n3346), .Y(n3345) );
  OR2X4 U3331 ( .A(n3277), .B(n3274), .Y(n3346) );
  OR2X4 U3332 ( .A(n3347), .B(n3348), .Y(n3274) );
  AND2X4 U3333 ( .A(n3349), .B(n3350), .Y(n3348) );
  AND2X4 U3334 ( .A(B[4]), .B(n3351), .Y(n3349) );
  OR2X4 U3335 ( .A(n131), .B(n3352), .Y(n3351) );
  OR2X4 U3336 ( .A(n3353), .B(n3354), .Y(n3352) );
  AND2X4 U3337 ( .A(n2233), .B(B[5]), .Y(n3354) );
  AND2X4 U3338 ( .A(A[2]), .B(n3355), .Y(n3353) );
  AND2X4 U3339 ( .A(n3356), .B(n3357), .Y(n3347) );
  OR2X4 U3340 ( .A(n3358), .B(n3359), .Y(n3356) );
  OR2X4 U3341 ( .A(n137), .B(n1241), .Y(n3359) );
  OR2X4 U3342 ( .A(n3360), .B(n3361), .Y(n3358) );
  AND2X4 U3343 ( .A(n141), .B(B[5]), .Y(n3361) );
  AND2X4 U3344 ( .A(n142), .B(n3355), .Y(n3360) );
  AND2X4 U3345 ( .A(A[3]), .B(B[3]), .Y(n3277) );
  INVX4 U3346 ( .A(n3278), .Y(n3279) );
  OR2X4 U3347 ( .A(n3362), .B(n3129), .Y(n3278) );
  INVX4 U3348 ( .A(B[3]), .Y(n3129) );
  AND2X4 U3349 ( .A(n3363), .B(n3364), .Y(n3362) );
  OR2X4 U3350 ( .A(n3365), .B(n1241), .Y(n3364) );
  AND2X4 U3351 ( .A(n2024), .B(n3366), .Y(n3365) );
  OR2X4 U3352 ( .A(n3246), .B(n1804), .Y(n3366) );
  OR2X4 U3353 ( .A(n3246), .B(n142), .Y(n3363) );
  INVX4 U3354 ( .A(n3252), .Y(n3246) );
  OR2X4 U3355 ( .A(n3367), .B(n3368), .Y(n3252) );
  AND2X4 U3356 ( .A(B[5]), .B(n3369), .Y(n3368) );
  OR2X4 U3357 ( .A(n3370), .B(n1207), .Y(n3369) );
  AND2X4 U3358 ( .A(A[0]), .B(n1241), .Y(n3370) );
  AND2X4 U3359 ( .A(B[4]), .B(n3371), .Y(n3367) );
  OR2X4 U3360 ( .A(n3372), .B(n1210), .Y(n3371) );
  AND2X4 U3361 ( .A(A[1]), .B(n3355), .Y(n3372) );
  OR2X4 U3362 ( .A(n3292), .B(n3289), .Y(n3344) );
  OR2X4 U3363 ( .A(n3373), .B(n3374), .Y(n3289) );
  OR2X4 U3364 ( .A(n3375), .B(n3376), .Y(n3374) );
  AND2X4 U3365 ( .A(n3377), .B(n3378), .Y(n3376) );
  INVX4 U3366 ( .A(n3379), .Y(n3378) );
  OR2X4 U3367 ( .A(n3380), .B(n3381), .Y(n3377) );
  AND2X4 U3368 ( .A(n3382), .B(n3383), .Y(n3381) );
  AND2X4 U3369 ( .A(n3384), .B(n3385), .Y(n3380) );
  AND2X4 U3370 ( .A(n3386), .B(n3379), .Y(n3375) );
  AND2X4 U3371 ( .A(n3385), .B(n3383), .Y(n3386) );
  INVX4 U3372 ( .A(n3382), .Y(n3385) );
  AND2X4 U3373 ( .A(n3387), .B(n3384), .Y(n3373) );
  AND2X4 U3374 ( .A(A[4]), .B(B[3]), .Y(n3292) );
  OR2X4 U3375 ( .A(n3307), .B(n3304), .Y(n3342) );
  OR2X4 U3376 ( .A(n3388), .B(n3389), .Y(n3304) );
  OR2X4 U3377 ( .A(n3390), .B(n3391), .Y(n3389) );
  AND2X4 U3378 ( .A(n3392), .B(n3393), .Y(n3391) );
  INVX4 U3379 ( .A(n3394), .Y(n3393) );
  AND2X4 U3380 ( .A(n3395), .B(n3396), .Y(n3392) );
  OR2X4 U3381 ( .A(n3397), .B(n3398), .Y(n3396) );
  OR2X4 U3382 ( .A(n3399), .B(n3400), .Y(n3395) );
  AND2X4 U3383 ( .A(n3401), .B(n3394), .Y(n3390) );
  AND2X4 U3384 ( .A(n3399), .B(n3400), .Y(n3401) );
  INVX4 U3385 ( .A(n3397), .Y(n3400) );
  INVX4 U3386 ( .A(n3398), .Y(n3399) );
  AND2X4 U3387 ( .A(n3402), .B(n3398), .Y(n3388) );
  AND2X4 U3388 ( .A(A[5]), .B(B[3]), .Y(n3307) );
  OR2X4 U3389 ( .A(n3322), .B(n3319), .Y(n3340) );
  OR2X4 U3390 ( .A(n3403), .B(n3404), .Y(n3319) );
  OR2X4 U3391 ( .A(n3405), .B(n3406), .Y(n3404) );
  AND2X4 U3392 ( .A(n3407), .B(n3408), .Y(n3406) );
  INVX4 U3393 ( .A(n3409), .Y(n3408) );
  AND2X4 U3394 ( .A(n3410), .B(n3411), .Y(n3407) );
  OR2X4 U3395 ( .A(n3412), .B(n3413), .Y(n3411) );
  OR2X4 U3396 ( .A(n3414), .B(n3415), .Y(n3410) );
  AND2X4 U3397 ( .A(n3416), .B(n3409), .Y(n3405) );
  AND2X4 U3398 ( .A(n3414), .B(n3415), .Y(n3416) );
  INVX4 U3399 ( .A(n3412), .Y(n3415) );
  INVX4 U3400 ( .A(n3413), .Y(n3414) );
  AND2X4 U3401 ( .A(n3417), .B(n3413), .Y(n3403) );
  AND2X4 U3402 ( .A(B[3]), .B(A[6]), .Y(n3322) );
  OR2X4 U3403 ( .A(n3418), .B(n3419), .Y(n2866) );
  AND2X4 U3404 ( .A(n3420), .B(n3421), .Y(n3419) );
  AND2X4 U3405 ( .A(n3422), .B(n2882), .Y(n3421) );
  OR2X4 U3406 ( .A(n3423), .B(n3424), .Y(n2882) );
  OR2X4 U3407 ( .A(n3425), .B(n3426), .Y(n3422) );
  INVX4 U3408 ( .A(n2881), .Y(n3420) );
  AND2X4 U3409 ( .A(n2881), .B(n3427), .Y(n3418) );
  OR2X4 U3410 ( .A(n3428), .B(n2880), .Y(n3427) );
  AND2X4 U3411 ( .A(n3424), .B(n3423), .Y(n2880) );
  AND2X4 U3412 ( .A(n3425), .B(n3426), .Y(n3428) );
  INVX4 U3413 ( .A(n3423), .Y(n3426) );
  AND2X4 U3414 ( .A(B[4]), .B(A[6]), .Y(n3423) );
  INVX4 U3415 ( .A(n3424), .Y(n3425) );
  OR2X4 U3416 ( .A(n3429), .B(n3417), .Y(n3424) );
  AND2X4 U3417 ( .A(n3409), .B(n3412), .Y(n3417) );
  AND2X4 U3418 ( .A(n3430), .B(n3413), .Y(n3429) );
  OR2X4 U3419 ( .A(n3431), .B(n3402), .Y(n3413) );
  AND2X4 U3420 ( .A(n3394), .B(n3397), .Y(n3402) );
  AND2X4 U3421 ( .A(n3432), .B(n3398), .Y(n3431) );
  OR2X4 U3422 ( .A(n3433), .B(n3387), .Y(n3398) );
  AND2X4 U3423 ( .A(n3379), .B(n3382), .Y(n3387) );
  AND2X4 U3424 ( .A(n3384), .B(n3434), .Y(n3433) );
  OR2X4 U3425 ( .A(n3382), .B(n3379), .Y(n3434) );
  OR2X4 U3426 ( .A(n3435), .B(n3436), .Y(n3379) );
  AND2X4 U3427 ( .A(n3437), .B(n3438), .Y(n3436) );
  AND2X4 U3428 ( .A(B[5]), .B(n3439), .Y(n3437) );
  OR2X4 U3429 ( .A(n131), .B(n3440), .Y(n3439) );
  OR2X4 U3430 ( .A(n3441), .B(n3442), .Y(n3440) );
  AND2X4 U3431 ( .A(n2233), .B(B[6]), .Y(n3442) );
  AND2X4 U3432 ( .A(A[2]), .B(n903), .Y(n3441) );
  AND2X4 U3433 ( .A(n3443), .B(n3444), .Y(n3435) );
  OR2X4 U3434 ( .A(n3445), .B(n3446), .Y(n3443) );
  OR2X4 U3435 ( .A(n137), .B(n3355), .Y(n3446) );
  OR2X4 U3436 ( .A(n3447), .B(n3448), .Y(n3445) );
  AND2X4 U3437 ( .A(n141), .B(B[6]), .Y(n3448) );
  AND2X4 U3438 ( .A(n142), .B(n903), .Y(n3447) );
  AND2X4 U3439 ( .A(A[3]), .B(B[4]), .Y(n3382) );
  INVX4 U3440 ( .A(n3383), .Y(n3384) );
  OR2X4 U3441 ( .A(n3449), .B(n1241), .Y(n3383) );
  INVX4 U3442 ( .A(B[4]), .Y(n1241) );
  AND2X4 U3443 ( .A(n3450), .B(n3451), .Y(n3449) );
  OR2X4 U3444 ( .A(n3452), .B(n3355), .Y(n3451) );
  AND2X4 U3445 ( .A(n2024), .B(n3453), .Y(n3452) );
  OR2X4 U3446 ( .A(n3350), .B(n1804), .Y(n3453) );
  OR2X4 U3447 ( .A(n3350), .B(n142), .Y(n3450) );
  INVX4 U3448 ( .A(n3357), .Y(n3350) );
  OR2X4 U3449 ( .A(n3454), .B(n3455), .Y(n3357) );
  AND2X4 U3450 ( .A(B[6]), .B(n3456), .Y(n3455) );
  OR2X4 U3451 ( .A(n3457), .B(n1207), .Y(n3456) );
  AND2X4 U3452 ( .A(A[0]), .B(n3355), .Y(n3457) );
  AND2X4 U3453 ( .A(B[5]), .B(n3458), .Y(n3454) );
  OR2X4 U3454 ( .A(n3459), .B(n1210), .Y(n3458) );
  AND2X4 U3455 ( .A(A[1]), .B(n903), .Y(n3459) );
  OR2X4 U3456 ( .A(n3397), .B(n3394), .Y(n3432) );
  OR2X4 U3457 ( .A(n3460), .B(n3461), .Y(n3394) );
  OR2X4 U3458 ( .A(n3462), .B(n3463), .Y(n3461) );
  AND2X4 U3459 ( .A(n3464), .B(n3465), .Y(n3463) );
  INVX4 U3460 ( .A(n3466), .Y(n3465) );
  OR2X4 U3461 ( .A(n3467), .B(n3468), .Y(n3464) );
  AND2X4 U3462 ( .A(n3469), .B(n3470), .Y(n3468) );
  AND2X4 U3463 ( .A(n3471), .B(n3472), .Y(n3467) );
  AND2X4 U3464 ( .A(n3473), .B(n3466), .Y(n3462) );
  AND2X4 U3465 ( .A(n3472), .B(n3470), .Y(n3473) );
  INVX4 U3466 ( .A(n3469), .Y(n3472) );
  AND2X4 U3467 ( .A(n3474), .B(n3471), .Y(n3460) );
  AND2X4 U3468 ( .A(A[4]), .B(B[4]), .Y(n3397) );
  OR2X4 U3469 ( .A(n3412), .B(n3409), .Y(n3430) );
  OR2X4 U3470 ( .A(n3475), .B(n3476), .Y(n3409) );
  OR2X4 U3471 ( .A(n3477), .B(n3478), .Y(n3476) );
  AND2X4 U3472 ( .A(n3479), .B(n3480), .Y(n3478) );
  INVX4 U3473 ( .A(n3481), .Y(n3480) );
  AND2X4 U3474 ( .A(n3482), .B(n3483), .Y(n3479) );
  OR2X4 U3475 ( .A(n3484), .B(n3485), .Y(n3483) );
  OR2X4 U3476 ( .A(n3486), .B(n3487), .Y(n3482) );
  AND2X4 U3477 ( .A(n3488), .B(n3481), .Y(n3477) );
  AND2X4 U3478 ( .A(n3486), .B(n3487), .Y(n3488) );
  INVX4 U3479 ( .A(n3484), .Y(n3487) );
  INVX4 U3480 ( .A(n3485), .Y(n3486) );
  AND2X4 U3481 ( .A(n3489), .B(n3485), .Y(n3475) );
  AND2X4 U3482 ( .A(B[4]), .B(A[5]), .Y(n3412) );
  OR2X4 U3483 ( .A(n3490), .B(n3491), .Y(n2881) );
  AND2X4 U3484 ( .A(n3492), .B(n3493), .Y(n3491) );
  AND2X4 U3485 ( .A(n3494), .B(n2897), .Y(n3493) );
  OR2X4 U3486 ( .A(n3495), .B(n3496), .Y(n2897) );
  OR2X4 U3487 ( .A(n3497), .B(n3498), .Y(n3494) );
  INVX4 U3488 ( .A(n2896), .Y(n3492) );
  AND2X4 U3489 ( .A(n2896), .B(n3499), .Y(n3490) );
  OR2X4 U3490 ( .A(n3500), .B(n2895), .Y(n3499) );
  AND2X4 U3491 ( .A(n3496), .B(n3495), .Y(n2895) );
  AND2X4 U3492 ( .A(n3497), .B(n3498), .Y(n3500) );
  INVX4 U3493 ( .A(n3495), .Y(n3498) );
  AND2X4 U3494 ( .A(B[5]), .B(A[5]), .Y(n3495) );
  INVX4 U3495 ( .A(n3496), .Y(n3497) );
  OR2X4 U3496 ( .A(n3501), .B(n3489), .Y(n3496) );
  AND2X4 U3497 ( .A(n3481), .B(n3484), .Y(n3489) );
  AND2X4 U3498 ( .A(n3502), .B(n3485), .Y(n3501) );
  OR2X4 U3499 ( .A(n3503), .B(n3474), .Y(n3485) );
  AND2X4 U3500 ( .A(n3466), .B(n3469), .Y(n3474) );
  AND2X4 U3501 ( .A(n3471), .B(n3504), .Y(n3503) );
  OR2X4 U3502 ( .A(n3469), .B(n3466), .Y(n3504) );
  OR2X4 U3503 ( .A(n3505), .B(n3506), .Y(n3466) );
  AND2X4 U3504 ( .A(n3507), .B(n3508), .Y(n3506) );
  AND2X4 U3505 ( .A(B[6]), .B(n3509), .Y(n3507) );
  OR2X4 U3506 ( .A(n131), .B(n3510), .Y(n3509) );
  OR2X4 U3507 ( .A(n3511), .B(n3512), .Y(n3510) );
  AND2X4 U3508 ( .A(n2233), .B(B[7]), .Y(n3512) );
  AND2X4 U3509 ( .A(A[2]), .B(n3513), .Y(n3511) );
  AND2X4 U3510 ( .A(n3514), .B(n3515), .Y(n3505) );
  OR2X4 U3511 ( .A(n3516), .B(n3517), .Y(n3514) );
  OR2X4 U3512 ( .A(n137), .B(n903), .Y(n3517) );
  OR2X4 U3513 ( .A(n3518), .B(n3519), .Y(n3516) );
  AND2X4 U3514 ( .A(n141), .B(B[7]), .Y(n3519) );
  AND2X4 U3515 ( .A(n142), .B(n3513), .Y(n3518) );
  AND2X4 U3516 ( .A(A[3]), .B(B[5]), .Y(n3469) );
  INVX4 U3517 ( .A(n3470), .Y(n3471) );
  OR2X4 U3518 ( .A(n3520), .B(n3355), .Y(n3470) );
  INVX4 U3519 ( .A(B[5]), .Y(n3355) );
  AND2X4 U3520 ( .A(n3521), .B(n3522), .Y(n3520) );
  OR2X4 U3521 ( .A(n3523), .B(n903), .Y(n3522) );
  AND2X4 U3522 ( .A(n2024), .B(n3524), .Y(n3523) );
  OR2X4 U3523 ( .A(n3438), .B(n1804), .Y(n3524) );
  OR2X4 U3524 ( .A(n3438), .B(n142), .Y(n3521) );
  INVX4 U3525 ( .A(n3444), .Y(n3438) );
  OR2X4 U3526 ( .A(n3525), .B(n3526), .Y(n3444) );
  AND2X4 U3527 ( .A(B[7]), .B(n3527), .Y(n3526) );
  OR2X4 U3528 ( .A(n3528), .B(n1207), .Y(n3527) );
  AND2X4 U3529 ( .A(A[0]), .B(n903), .Y(n3528) );
  AND2X4 U3530 ( .A(B[6]), .B(n3529), .Y(n3525) );
  OR2X4 U3531 ( .A(n3530), .B(n1210), .Y(n3529) );
  AND2X4 U3532 ( .A(A[1]), .B(n3513), .Y(n3530) );
  OR2X4 U3533 ( .A(n3484), .B(n3481), .Y(n3502) );
  OR2X4 U3534 ( .A(n3531), .B(n3532), .Y(n3481) );
  OR2X4 U3535 ( .A(n3533), .B(n3534), .Y(n3532) );
  AND2X4 U3536 ( .A(n3535), .B(n3536), .Y(n3534) );
  INVX4 U3537 ( .A(n3537), .Y(n3536) );
  OR2X4 U3538 ( .A(n3538), .B(n3539), .Y(n3535) );
  AND2X4 U3539 ( .A(n3540), .B(n3541), .Y(n3539) );
  AND2X4 U3540 ( .A(n3542), .B(n3543), .Y(n3538) );
  AND2X4 U3541 ( .A(n3544), .B(n3537), .Y(n3533) );
  AND2X4 U3542 ( .A(n3543), .B(n3541), .Y(n3544) );
  INVX4 U3543 ( .A(n3540), .Y(n3543) );
  AND2X4 U3544 ( .A(n3545), .B(n3542), .Y(n3531) );
  AND2X4 U3545 ( .A(B[5]), .B(A[4]), .Y(n3484) );
  OR2X4 U3546 ( .A(n3546), .B(n3547), .Y(n2896) );
  AND2X4 U3547 ( .A(n3548), .B(n3549), .Y(n3547) );
  AND2X4 U3548 ( .A(n3550), .B(n2912), .Y(n3549) );
  OR2X4 U3549 ( .A(n3551), .B(n3552), .Y(n2912) );
  OR2X4 U3550 ( .A(n3553), .B(n3554), .Y(n3550) );
  INVX4 U3551 ( .A(n2911), .Y(n3548) );
  AND2X4 U3552 ( .A(n2911), .B(n3555), .Y(n3546) );
  OR2X4 U3553 ( .A(n3556), .B(n2910), .Y(n3555) );
  AND2X4 U3554 ( .A(n3552), .B(n3551), .Y(n2910) );
  AND2X4 U3555 ( .A(n3553), .B(n3554), .Y(n3556) );
  INVX4 U3556 ( .A(n3551), .Y(n3554) );
  AND2X4 U3557 ( .A(B[6]), .B(A[4]), .Y(n3551) );
  INVX4 U3558 ( .A(n3552), .Y(n3553) );
  OR2X4 U3559 ( .A(n3557), .B(n3545), .Y(n3552) );
  AND2X4 U3560 ( .A(n3537), .B(n3540), .Y(n3545) );
  AND2X4 U3561 ( .A(n3542), .B(n3558), .Y(n3557) );
  OR2X4 U3562 ( .A(n3540), .B(n3537), .Y(n3558) );
  OR2X4 U3563 ( .A(n3559), .B(n3560), .Y(n3537) );
  AND2X4 U3564 ( .A(n3561), .B(n3562), .Y(n3560) );
  AND2X4 U3565 ( .A(B[7]), .B(n3563), .Y(n3561) );
  OR2X4 U3566 ( .A(n131), .B(n3564), .Y(n3563) );
  OR2X4 U3567 ( .A(n3565), .B(n3566), .Y(n3564) );
  AND2X4 U3568 ( .A(n2233), .B(B[8]), .Y(n3566) );
  AND2X4 U3569 ( .A(A[2]), .B(n633), .Y(n3565) );
  AND2X4 U3570 ( .A(n3567), .B(n3568), .Y(n3559) );
  OR2X4 U3571 ( .A(n3569), .B(n3570), .Y(n3567) );
  OR2X4 U3572 ( .A(n137), .B(n3513), .Y(n3570) );
  OR2X4 U3573 ( .A(n3571), .B(n3572), .Y(n3569) );
  AND2X4 U3574 ( .A(n141), .B(B[8]), .Y(n3572) );
  AND2X4 U3575 ( .A(n142), .B(n633), .Y(n3571) );
  AND2X4 U3576 ( .A(B[6]), .B(A[3]), .Y(n3540) );
  INVX4 U3577 ( .A(n3541), .Y(n3542) );
  OR2X4 U3578 ( .A(n3573), .B(n903), .Y(n3541) );
  INVX4 U3579 ( .A(B[6]), .Y(n903) );
  AND2X4 U3580 ( .A(n3574), .B(n3575), .Y(n3573) );
  OR2X4 U3581 ( .A(n3576), .B(n3513), .Y(n3575) );
  AND2X4 U3582 ( .A(n2024), .B(n3577), .Y(n3576) );
  OR2X4 U3583 ( .A(n3508), .B(n1804), .Y(n3577) );
  OR2X4 U3584 ( .A(n3508), .B(n142), .Y(n3574) );
  INVX4 U3585 ( .A(n3515), .Y(n3508) );
  OR2X4 U3586 ( .A(n3578), .B(n3579), .Y(n3515) );
  AND2X4 U3587 ( .A(B[8]), .B(n3580), .Y(n3579) );
  OR2X4 U3588 ( .A(n3581), .B(n1207), .Y(n3580) );
  AND2X4 U3589 ( .A(A[0]), .B(n3513), .Y(n3581) );
  AND2X4 U3590 ( .A(B[7]), .B(n3582), .Y(n3578) );
  OR2X4 U3591 ( .A(n3583), .B(n1210), .Y(n3582) );
  AND2X4 U3592 ( .A(A[1]), .B(n633), .Y(n3583) );
  OR2X4 U3593 ( .A(n3584), .B(n3585), .Y(n2911) );
  AND2X4 U3594 ( .A(n3586), .B(n3587), .Y(n3585) );
  INVX4 U3595 ( .A(n2926), .Y(n3587) );
  OR2X4 U3596 ( .A(n3588), .B(n3589), .Y(n3586) );
  AND2X4 U3597 ( .A(n2928), .B(n3590), .Y(n3589) );
  AND2X4 U3598 ( .A(n2929), .B(n3591), .Y(n3588) );
  AND2X4 U3599 ( .A(n2926), .B(n3592), .Y(n3584) );
  OR2X4 U3600 ( .A(n3593), .B(n2925), .Y(n3592) );
  AND2X4 U3601 ( .A(n2928), .B(n2929), .Y(n2925) );
  INVX4 U3602 ( .A(n3590), .Y(n2929) );
  AND2X4 U3603 ( .A(n3591), .B(n3590), .Y(n3593) );
  OR2X4 U3604 ( .A(n3594), .B(n3513), .Y(n3590) );
  INVX4 U3605 ( .A(B[7]), .Y(n3513) );
  AND2X4 U3606 ( .A(n3595), .B(n3596), .Y(n3594) );
  OR2X4 U3607 ( .A(n3597), .B(n633), .Y(n3596) );
  AND2X4 U3608 ( .A(n2024), .B(n3598), .Y(n3597) );
  OR2X4 U3609 ( .A(n3562), .B(n1804), .Y(n3598) );
  INVX4 U3610 ( .A(n141), .Y(n2024) );
  OR2X4 U3611 ( .A(n3562), .B(n142), .Y(n3595) );
  INVX4 U3612 ( .A(n3568), .Y(n3562) );
  OR2X4 U3613 ( .A(n3599), .B(n3600), .Y(n3568) );
  AND2X4 U3614 ( .A(B[9]), .B(n3601), .Y(n3600) );
  OR2X4 U3615 ( .A(n3602), .B(n1207), .Y(n3601) );
  AND2X4 U3616 ( .A(A[0]), .B(n633), .Y(n3602) );
  AND2X4 U3617 ( .A(B[8]), .B(n3603), .Y(n3599) );
  OR2X4 U3618 ( .A(n3604), .B(n1210), .Y(n3603) );
  AND2X4 U3619 ( .A(A[1]), .B(n2783), .Y(n3604) );
  INVX4 U3620 ( .A(n2928), .Y(n3591) );
  AND2X4 U3621 ( .A(B[7]), .B(A[3]), .Y(n2928) );
  OR2X4 U3622 ( .A(n3605), .B(n3606), .Y(n2926) );
  AND2X4 U3623 ( .A(n3607), .B(n2945), .Y(n3606) );
  INVX4 U3624 ( .A(n3608), .Y(n2945) );
  AND2X4 U3625 ( .A(B[8]), .B(n3609), .Y(n3607) );
  OR2X4 U3626 ( .A(n131), .B(n3610), .Y(n3609) );
  OR2X4 U3627 ( .A(n3611), .B(n3612), .Y(n3610) );
  AND2X4 U3628 ( .A(n2233), .B(B[9]), .Y(n3612) );
  AND2X4 U3629 ( .A(n142), .B(n3613), .Y(n2233) );
  AND2X4 U3630 ( .A(A[2]), .B(n2783), .Y(n3611) );
  AND2X4 U3631 ( .A(n1804), .B(A[2]), .Y(n131) );
  AND2X4 U3632 ( .A(n3614), .B(n3608), .Y(n3605) );
  OR2X4 U3633 ( .A(n3615), .B(n3616), .Y(n3608) );
  AND2X4 U3634 ( .A(B[9]), .B(n3617), .Y(n3616) );
  OR2X4 U3635 ( .A(n3618), .B(n1210), .Y(n3617) );
  NOR2X4 U3636 ( .A(A[0]), .B(n1806), .Y(n1210) );
  AND2X4 U3637 ( .A(A[1]), .B(n423), .Y(n3618) );
  INVX4 U3638 ( .A(B[10]), .Y(n423) );
  AND2X4 U3639 ( .A(B[10]), .B(n3619), .Y(n3615) );
  OR2X4 U3640 ( .A(n3620), .B(n1207), .Y(n3619) );
  AND2X4 U3641 ( .A(n1806), .B(A[0]), .Y(n1207) );
  INVX4 U3642 ( .A(A[1]), .Y(n1806) );
  AND2X4 U3643 ( .A(A[0]), .B(n2783), .Y(n3620) );
  OR2X4 U3644 ( .A(n3621), .B(n3622), .Y(n3614) );
  OR2X4 U3645 ( .A(n137), .B(n633), .Y(n3622) );
  INVX4 U3646 ( .A(B[8]), .Y(n633) );
  AND2X4 U3647 ( .A(n142), .B(n1804), .Y(n137) );
  INVX4 U3648 ( .A(n3613), .Y(n1804) );
  OR2X4 U3649 ( .A(n3623), .B(n3624), .Y(n3621) );
  AND2X4 U3650 ( .A(n141), .B(B[9]), .Y(n3624) );
  AND2X4 U3651 ( .A(n3613), .B(A[2]), .Y(n141) );
  AND2X4 U3652 ( .A(A[0]), .B(A[1]), .Y(n3613) );
  AND2X4 U3653 ( .A(n142), .B(n2783), .Y(n3623) );
  INVX4 U3654 ( .A(B[9]), .Y(n2783) );
  INVX4 U3655 ( .A(A[2]), .Y(n142) );
  AND2X4 U3656 ( .A(A[0]), .B(B[0]), .Y(Y[0]) );
endmodule

